magic
tech scmos
timestamp 1764437107
<< nwell >>
rect -130 1777 -97 1870
rect -78 1791 -54 1843
rect -18 1791 8 1843
rect 42 1777 66 1829
rect 672 1765 705 1858
rect 724 1779 748 1831
rect 784 1779 810 1831
rect 844 1765 868 1817
rect 250 1704 302 1736
rect 94 1639 146 1671
rect 416 1667 468 1699
rect -200 1527 -167 1620
rect 250 1618 302 1650
rect -148 1541 -124 1593
rect -88 1541 -62 1593
rect -28 1527 -4 1579
rect 609 1567 633 1623
rect 1758 1618 1810 1650
rect 2170 1626 2203 1719
rect 2222 1640 2246 1692
rect 2282 1640 2308 1692
rect 2342 1626 2366 1678
rect 222 1529 274 1561
rect 1602 1553 1654 1585
rect 1924 1581 1976 1613
rect 1758 1532 1810 1564
rect -525 1300 -492 1393
rect -473 1314 -449 1366
rect -413 1314 -387 1366
rect -353 1300 -329 1352
rect -168 1303 -135 1396
rect -116 1317 -92 1369
rect -56 1317 -30 1369
rect 4 1303 28 1355
rect 257 1353 309 1385
rect 101 1288 153 1320
rect 423 1316 475 1348
rect 1758 1343 1810 1375
rect 2174 1366 2207 1459
rect 2226 1380 2250 1432
rect 2286 1380 2312 1432
rect 2346 1366 2370 1418
rect 257 1267 309 1299
rect 965 1283 1017 1315
rect 1602 1278 1654 1310
rect 1924 1306 1976 1338
rect 612 1216 636 1272
rect 1758 1257 1810 1289
rect 1189 1218 1241 1250
rect 229 1178 281 1210
rect 1760 1149 1812 1181
rect -549 986 -516 1079
rect -497 1000 -473 1052
rect -437 1000 -411 1052
rect -377 986 -353 1038
rect -218 996 -185 1089
rect 959 1080 1011 1108
rect 1604 1084 1656 1116
rect 1926 1112 1978 1144
rect 2182 1142 2215 1235
rect 2234 1156 2258 1208
rect 2294 1156 2320 1208
rect 2354 1142 2378 1194
rect 958 1068 1011 1080
rect -166 1010 -142 1062
rect -106 1010 -80 1062
rect -46 996 -22 1048
rect 227 1012 279 1044
rect 1148 1039 1200 1067
rect 1760 1063 1812 1095
rect 1147 1027 1200 1039
rect 71 947 123 979
rect 393 975 445 1007
rect 968 992 1020 1024
rect 227 926 279 958
rect 1767 948 1819 980
rect 591 875 615 931
rect 945 894 997 942
rect 199 837 251 869
rect 1164 845 1216 893
rect 1611 883 1663 915
rect 1933 911 1985 943
rect 2175 922 2208 1015
rect 2227 936 2251 988
rect 2287 936 2313 988
rect 2347 922 2371 974
rect 1767 862 1819 894
rect 955 817 1007 845
rect 954 805 1007 817
rect -508 644 -475 737
rect -456 658 -432 710
rect -396 658 -370 710
rect -336 644 -312 696
rect -199 648 -166 741
rect 964 740 1016 772
rect -147 662 -123 714
rect -87 662 -61 714
rect -27 648 -3 700
rect 226 670 278 702
rect 70 605 122 637
rect 392 633 444 665
rect 226 584 278 616
rect 585 533 609 589
rect 198 495 250 527
rect -589 313 -556 406
rect -537 327 -513 379
rect -477 327 -451 379
rect -417 313 -393 365
rect -251 313 -218 406
rect 220 388 272 420
rect -199 327 -175 379
rect -139 327 -113 379
rect -79 313 -55 365
rect 64 323 116 355
rect 386 351 438 383
rect 913 380 965 436
rect 220 302 272 334
rect 1197 295 1249 351
rect 192 213 244 245
rect 935 227 987 275
rect 1618 261 1651 354
rect 1670 275 1694 327
rect 1730 275 1756 327
rect 1790 261 1814 313
rect 948 103 1000 131
rect 947 91 1000 103
rect 968 9 1020 41
<< ntransistor >>
rect -119 1728 -117 1748
rect -67 1742 -65 1782
rect -59 1742 -57 1782
rect -7 1742 -5 1782
rect 1 1742 3 1782
rect 53 1749 55 1769
rect 311 1723 351 1725
rect 311 1715 351 1717
rect 683 1716 685 1736
rect 735 1730 737 1770
rect 743 1730 745 1770
rect 795 1730 797 1770
rect 803 1730 805 1770
rect 855 1737 857 1757
rect 477 1686 517 1688
rect 477 1678 517 1680
rect 155 1658 195 1660
rect 155 1650 195 1652
rect 311 1637 351 1639
rect 1819 1637 1859 1639
rect 311 1629 351 1631
rect 1819 1629 1859 1631
rect 1985 1600 2025 1602
rect 1985 1592 2025 1594
rect 2181 1577 2183 1597
rect 2233 1591 2235 1631
rect 2241 1591 2243 1631
rect 2293 1591 2295 1631
rect 2301 1591 2303 1631
rect 2353 1598 2355 1618
rect 1663 1572 1703 1574
rect 1663 1564 1703 1566
rect 283 1548 323 1550
rect 283 1540 323 1542
rect 620 1539 622 1559
rect 1819 1551 1859 1553
rect 1819 1543 1859 1545
rect -189 1478 -187 1498
rect -137 1492 -135 1532
rect -129 1492 -127 1532
rect -77 1492 -75 1532
rect -69 1492 -67 1532
rect -17 1499 -15 1519
rect 318 1372 358 1374
rect 318 1364 358 1366
rect 1819 1362 1859 1364
rect 1819 1354 1859 1356
rect -514 1251 -512 1271
rect -462 1265 -460 1305
rect -454 1265 -452 1305
rect -402 1265 -400 1305
rect -394 1265 -392 1305
rect -342 1272 -340 1292
rect 484 1335 524 1337
rect 484 1327 524 1329
rect 1985 1325 2025 1327
rect 1985 1317 2025 1319
rect 2185 1317 2187 1337
rect 2237 1331 2239 1371
rect 2245 1331 2247 1371
rect 2297 1331 2299 1371
rect 2305 1331 2307 1371
rect 2357 1338 2359 1358
rect -157 1254 -155 1274
rect -105 1268 -103 1308
rect -97 1268 -95 1308
rect -45 1268 -43 1308
rect -37 1268 -35 1308
rect 162 1307 202 1309
rect 1026 1302 1066 1304
rect 162 1299 202 1301
rect 15 1275 17 1295
rect 1663 1297 1703 1299
rect 1026 1294 1066 1296
rect 1663 1289 1703 1291
rect 318 1286 358 1288
rect 318 1278 358 1280
rect 1819 1276 1859 1278
rect 1819 1268 1859 1270
rect 1250 1237 1290 1239
rect 1250 1229 1290 1231
rect 290 1197 330 1199
rect 290 1189 330 1191
rect 623 1188 625 1208
rect 1821 1168 1861 1170
rect 1821 1160 1861 1162
rect 1987 1131 2027 1133
rect 1987 1123 2027 1125
rect 1665 1103 1705 1105
rect 1023 1095 1083 1097
rect 1665 1095 1705 1097
rect 2193 1093 2195 1113
rect 2245 1107 2247 1147
rect 2253 1107 2255 1147
rect 2305 1107 2307 1147
rect 2313 1107 2315 1147
rect 2365 1114 2367 1134
rect 1023 1087 1083 1089
rect 1821 1082 1861 1084
rect 1023 1079 1083 1081
rect 1821 1074 1861 1076
rect 1212 1054 1272 1056
rect 1212 1046 1272 1048
rect -538 937 -536 957
rect -486 951 -484 991
rect -478 951 -476 991
rect -426 951 -424 991
rect -418 951 -416 991
rect -366 958 -364 978
rect 1212 1038 1272 1040
rect 288 1031 328 1033
rect 288 1023 328 1025
rect 1029 1011 1069 1013
rect 1029 1003 1069 1005
rect -207 947 -205 967
rect -155 961 -153 1001
rect -147 961 -145 1001
rect -95 961 -93 1001
rect -87 961 -85 1001
rect 454 994 494 996
rect -35 968 -33 988
rect 454 986 494 988
rect 132 966 172 968
rect 1828 967 1868 969
rect 132 958 172 960
rect 1828 959 1868 961
rect 288 945 328 947
rect 288 937 328 939
rect 1015 929 1095 931
rect 1994 930 2034 932
rect 1015 921 1095 923
rect 1994 922 2034 924
rect 1015 913 1095 915
rect 1015 905 1095 907
rect 1672 902 1712 904
rect 1672 894 1712 896
rect 1234 880 1314 882
rect 1828 881 1868 883
rect 1234 872 1314 874
rect 1828 873 1868 875
rect 2186 873 2188 893
rect 2238 887 2240 927
rect 2246 887 2248 927
rect 2298 887 2300 927
rect 2306 887 2308 927
rect 2358 894 2360 914
rect 260 856 300 858
rect 260 848 300 850
rect 602 847 604 867
rect 1234 864 1314 866
rect 1234 856 1314 858
rect 1019 832 1079 834
rect 1019 824 1079 826
rect 1019 816 1079 818
rect 1025 759 1065 761
rect 1025 751 1065 753
rect -497 595 -495 615
rect -445 609 -443 649
rect -437 609 -435 649
rect -385 609 -383 649
rect -377 609 -375 649
rect -325 616 -323 636
rect 287 689 327 691
rect 287 681 327 683
rect -188 599 -186 619
rect -136 613 -134 653
rect -128 613 -126 653
rect -76 613 -74 653
rect -68 613 -66 653
rect 453 652 493 654
rect 453 644 493 646
rect -16 620 -14 640
rect 131 624 171 626
rect 131 616 171 618
rect 287 603 327 605
rect 287 595 327 597
rect 259 514 299 516
rect 259 506 299 508
rect 596 505 598 525
rect 983 423 1063 425
rect 983 415 1063 417
rect 281 407 321 409
rect 983 407 1063 409
rect 281 399 321 401
rect 983 399 1063 401
rect 983 391 1063 393
rect 447 370 487 372
rect 447 362 487 364
rect -578 264 -576 284
rect -526 278 -524 318
rect -518 278 -516 318
rect -466 278 -464 318
rect -458 278 -456 318
rect -406 285 -404 305
rect 125 342 165 344
rect 1267 338 1347 340
rect 125 334 165 336
rect 1267 330 1347 332
rect 281 321 321 323
rect 1267 322 1347 324
rect -240 264 -238 284
rect -188 278 -186 318
rect -180 278 -178 318
rect -128 278 -126 318
rect -120 278 -118 318
rect 281 313 321 315
rect 1267 314 1347 316
rect 1267 306 1347 308
rect -68 285 -66 305
rect 1005 262 1085 264
rect 1005 254 1085 256
rect 1005 246 1085 248
rect 1005 238 1085 240
rect 253 232 293 234
rect 253 224 293 226
rect 1629 212 1631 232
rect 1681 226 1683 266
rect 1689 226 1691 266
rect 1741 226 1743 266
rect 1749 226 1751 266
rect 1801 233 1803 253
rect 1012 118 1072 120
rect 1012 110 1072 112
rect 1012 102 1072 104
rect 1029 28 1069 30
rect 1029 20 1069 22
<< ptransistor >>
rect -119 1784 -117 1864
rect -111 1784 -109 1864
rect -67 1797 -65 1837
rect -7 1797 -5 1837
rect 53 1783 55 1823
rect 683 1772 685 1852
rect 691 1772 693 1852
rect 735 1785 737 1825
rect 795 1785 797 1825
rect 855 1771 857 1811
rect 256 1723 296 1725
rect 256 1715 296 1717
rect 422 1686 462 1688
rect 422 1678 462 1680
rect 100 1658 140 1660
rect 100 1650 140 1652
rect 256 1637 296 1639
rect 1764 1637 1804 1639
rect 256 1629 296 1631
rect 2181 1633 2183 1713
rect 2189 1633 2191 1713
rect 2233 1646 2235 1686
rect 2293 1646 2295 1686
rect 1764 1629 1804 1631
rect -189 1534 -187 1614
rect -181 1534 -179 1614
rect -137 1547 -135 1587
rect -77 1547 -75 1587
rect 620 1573 622 1613
rect 1930 1600 1970 1602
rect 2353 1632 2355 1672
rect 1930 1592 1970 1594
rect -17 1533 -15 1573
rect 1608 1572 1648 1574
rect 1608 1564 1648 1566
rect 228 1548 268 1550
rect 228 1540 268 1542
rect 1764 1551 1804 1553
rect 1764 1543 1804 1545
rect -514 1307 -512 1387
rect -506 1307 -504 1387
rect -462 1320 -460 1360
rect -402 1320 -400 1360
rect -342 1306 -340 1346
rect -157 1310 -155 1390
rect -149 1310 -147 1390
rect 263 1372 303 1374
rect 2185 1373 2187 1453
rect 2193 1373 2195 1453
rect 2237 1386 2239 1426
rect 2297 1386 2299 1426
rect 263 1364 303 1366
rect -105 1323 -103 1363
rect -45 1323 -43 1363
rect 1764 1362 1804 1364
rect 1764 1354 1804 1356
rect 15 1309 17 1349
rect 2357 1372 2359 1412
rect 429 1335 469 1337
rect 429 1327 469 1329
rect 1930 1325 1970 1327
rect 1930 1317 1970 1319
rect 107 1307 147 1309
rect 971 1302 1011 1304
rect 107 1299 147 1301
rect 1608 1297 1648 1299
rect 971 1294 1011 1296
rect 1608 1289 1648 1291
rect 263 1286 303 1288
rect 263 1278 303 1280
rect 1764 1276 1804 1278
rect 1764 1268 1804 1270
rect 623 1222 625 1262
rect 1195 1237 1235 1239
rect 1195 1229 1235 1231
rect 235 1197 275 1199
rect 235 1189 275 1191
rect 1766 1168 1806 1170
rect 1766 1160 1806 1162
rect 2193 1149 2195 1229
rect 2201 1149 2203 1229
rect 2245 1162 2247 1202
rect 2305 1162 2307 1202
rect 1932 1131 1972 1133
rect 1932 1123 1972 1125
rect 2365 1148 2367 1188
rect 1610 1103 1650 1105
rect 965 1095 1005 1097
rect 1610 1095 1650 1097
rect 965 1087 1005 1089
rect -538 993 -536 1073
rect -530 993 -528 1073
rect -486 1006 -484 1046
rect -426 1006 -424 1046
rect -366 992 -364 1032
rect -207 1003 -205 1083
rect -199 1003 -197 1083
rect 1766 1082 1806 1084
rect 965 1079 1005 1081
rect 1766 1074 1806 1076
rect -155 1016 -153 1056
rect -95 1016 -93 1056
rect 1154 1054 1194 1056
rect 1154 1046 1194 1048
rect -35 1002 -33 1042
rect 1154 1038 1194 1040
rect 233 1031 273 1033
rect 233 1023 273 1025
rect 974 1011 1014 1013
rect 974 1003 1014 1005
rect 399 994 439 996
rect 399 986 439 988
rect 77 966 117 968
rect 1773 967 1813 969
rect 77 958 117 960
rect 1773 959 1813 961
rect 233 945 273 947
rect 233 937 273 939
rect 951 929 991 931
rect 1939 930 1979 932
rect 602 881 604 921
rect 951 921 991 923
rect 2186 929 2188 1009
rect 2194 929 2196 1009
rect 2238 942 2240 982
rect 2298 942 2300 982
rect 1939 922 1979 924
rect 951 913 991 915
rect 951 905 991 907
rect 1617 902 1657 904
rect 1617 894 1657 896
rect 2358 928 2360 968
rect 1170 880 1210 882
rect 1773 881 1813 883
rect 1170 872 1210 874
rect 1773 873 1813 875
rect 205 856 245 858
rect 205 848 245 850
rect 1170 864 1210 866
rect 1170 856 1210 858
rect 961 832 1001 834
rect 961 824 1001 826
rect 961 816 1001 818
rect 970 759 1010 761
rect 970 751 1010 753
rect -497 651 -495 731
rect -489 651 -487 731
rect -445 664 -443 704
rect -385 664 -383 704
rect -325 650 -323 690
rect -188 655 -186 735
rect -180 655 -178 735
rect -136 668 -134 708
rect -76 668 -74 708
rect -16 654 -14 694
rect 232 689 272 691
rect 232 681 272 683
rect 398 652 438 654
rect 398 644 438 646
rect 76 624 116 626
rect 76 616 116 618
rect 232 603 272 605
rect 232 595 272 597
rect 596 539 598 579
rect 204 514 244 516
rect 204 506 244 508
rect 919 423 959 425
rect 919 415 959 417
rect 226 407 266 409
rect -578 320 -576 400
rect -570 320 -568 400
rect -526 333 -524 373
rect -466 333 -464 373
rect -406 319 -404 359
rect -240 320 -238 400
rect -232 320 -230 400
rect 919 407 959 409
rect 226 399 266 401
rect 919 399 959 401
rect 919 391 959 393
rect -188 333 -186 373
rect -128 333 -126 373
rect 392 370 432 372
rect 392 362 432 364
rect -68 319 -66 359
rect 70 342 110 344
rect 1203 338 1243 340
rect 70 334 110 336
rect 1203 330 1243 332
rect 226 321 266 323
rect 1203 322 1243 324
rect 226 313 266 315
rect 1203 314 1243 316
rect 1203 306 1243 308
rect 1629 268 1631 348
rect 1637 268 1639 348
rect 1681 281 1683 321
rect 1741 281 1743 321
rect 941 262 981 264
rect 941 254 981 256
rect 941 246 981 248
rect 941 238 981 240
rect 198 232 238 234
rect 1801 267 1803 307
rect 198 224 238 226
rect 954 118 994 120
rect 954 110 994 112
rect 954 102 994 104
rect 974 28 1014 30
rect 974 20 1014 22
<< ndiffusion >>
rect -120 1728 -119 1748
rect -117 1728 -116 1748
rect -68 1742 -67 1782
rect -65 1742 -64 1782
rect -60 1742 -59 1782
rect -57 1742 -56 1782
rect -8 1742 -7 1782
rect -5 1742 -4 1782
rect 0 1742 1 1782
rect 3 1742 4 1782
rect 52 1749 53 1769
rect 55 1749 56 1769
rect 311 1725 351 1726
rect 311 1722 351 1723
rect 311 1717 351 1718
rect 682 1716 683 1736
rect 685 1716 686 1736
rect 734 1730 735 1770
rect 737 1730 738 1770
rect 742 1730 743 1770
rect 745 1730 746 1770
rect 794 1730 795 1770
rect 797 1730 798 1770
rect 802 1730 803 1770
rect 805 1730 806 1770
rect 854 1737 855 1757
rect 857 1737 858 1757
rect 311 1714 351 1715
rect 477 1688 517 1689
rect 477 1685 517 1686
rect 477 1680 517 1681
rect 477 1677 517 1678
rect 155 1660 195 1661
rect 155 1657 195 1658
rect 155 1652 195 1653
rect 155 1649 195 1650
rect 311 1639 351 1640
rect 311 1636 351 1637
rect 1819 1639 1859 1640
rect 311 1631 351 1632
rect 311 1628 351 1629
rect 1819 1636 1859 1637
rect 1819 1631 1859 1632
rect 1819 1628 1859 1629
rect 1985 1602 2025 1603
rect 1985 1599 2025 1600
rect 1985 1594 2025 1595
rect 1985 1591 2025 1592
rect 2180 1577 2181 1597
rect 2183 1577 2184 1597
rect 2232 1591 2233 1631
rect 2235 1591 2236 1631
rect 2240 1591 2241 1631
rect 2243 1591 2244 1631
rect 2292 1591 2293 1631
rect 2295 1591 2296 1631
rect 2300 1591 2301 1631
rect 2303 1591 2304 1631
rect 2352 1598 2353 1618
rect 2355 1598 2356 1618
rect 1663 1574 1703 1575
rect 1663 1571 1703 1572
rect 1663 1566 1703 1567
rect 1663 1563 1703 1564
rect 283 1550 323 1551
rect 283 1547 323 1548
rect 283 1542 323 1543
rect 283 1539 323 1540
rect 619 1539 620 1559
rect 622 1539 623 1559
rect 1819 1553 1859 1554
rect 1819 1550 1859 1551
rect 1819 1545 1859 1546
rect 1819 1542 1859 1543
rect -190 1478 -189 1498
rect -187 1478 -186 1498
rect -138 1492 -137 1532
rect -135 1492 -134 1532
rect -130 1492 -129 1532
rect -127 1492 -126 1532
rect -78 1492 -77 1532
rect -75 1492 -74 1532
rect -70 1492 -69 1532
rect -67 1492 -66 1532
rect -18 1499 -17 1519
rect -15 1499 -14 1519
rect 318 1374 358 1375
rect 318 1371 358 1372
rect 318 1366 358 1367
rect 318 1363 358 1364
rect 1819 1364 1859 1365
rect 1819 1361 1859 1362
rect 1819 1356 1859 1357
rect 1819 1353 1859 1354
rect -515 1251 -514 1271
rect -512 1251 -511 1271
rect -463 1265 -462 1305
rect -460 1265 -459 1305
rect -455 1265 -454 1305
rect -452 1265 -451 1305
rect -403 1265 -402 1305
rect -400 1265 -399 1305
rect -395 1265 -394 1305
rect -392 1265 -391 1305
rect -343 1272 -342 1292
rect -340 1272 -339 1292
rect 484 1337 524 1338
rect 484 1334 524 1335
rect 484 1329 524 1330
rect 484 1326 524 1327
rect 1985 1327 2025 1328
rect 1985 1324 2025 1325
rect 1985 1319 2025 1320
rect 2184 1317 2185 1337
rect 2187 1317 2188 1337
rect 2236 1331 2237 1371
rect 2239 1331 2240 1371
rect 2244 1331 2245 1371
rect 2247 1331 2248 1371
rect 2296 1331 2297 1371
rect 2299 1331 2300 1371
rect 2304 1331 2305 1371
rect 2307 1331 2308 1371
rect 2356 1338 2357 1358
rect 2359 1338 2360 1358
rect -158 1254 -157 1274
rect -155 1254 -154 1274
rect -106 1268 -105 1308
rect -103 1268 -102 1308
rect -98 1268 -97 1308
rect -95 1268 -94 1308
rect -46 1268 -45 1308
rect -43 1268 -42 1308
rect -38 1268 -37 1308
rect -35 1268 -34 1308
rect 1985 1316 2025 1317
rect 162 1309 202 1310
rect 162 1306 202 1307
rect 162 1301 202 1302
rect 1026 1304 1066 1305
rect 14 1275 15 1295
rect 17 1275 18 1295
rect 162 1298 202 1299
rect 1026 1301 1066 1302
rect 1026 1296 1066 1297
rect 1663 1299 1703 1300
rect 1026 1293 1066 1294
rect 318 1288 358 1289
rect 1663 1296 1703 1297
rect 1663 1291 1703 1292
rect 318 1285 358 1286
rect 1663 1288 1703 1289
rect 318 1280 358 1281
rect 318 1277 358 1278
rect 1819 1278 1859 1279
rect 1819 1275 1859 1276
rect 1819 1270 1859 1271
rect 1819 1267 1859 1268
rect 1250 1239 1290 1240
rect 1250 1236 1290 1237
rect 1250 1231 1290 1232
rect 1250 1228 1290 1229
rect 290 1199 330 1200
rect 290 1196 330 1197
rect 290 1191 330 1192
rect 290 1188 330 1189
rect 622 1188 623 1208
rect 625 1188 626 1208
rect 1821 1170 1861 1171
rect 1821 1167 1861 1168
rect 1821 1162 1861 1163
rect 1821 1159 1861 1160
rect 1987 1133 2027 1134
rect 1987 1130 2027 1131
rect 1987 1125 2027 1126
rect 1987 1122 2027 1123
rect 1665 1105 1705 1106
rect 1023 1097 1083 1098
rect 1023 1094 1083 1095
rect 1665 1102 1705 1103
rect 1665 1097 1705 1098
rect 1665 1094 1705 1095
rect 2192 1093 2193 1113
rect 2195 1093 2196 1113
rect 2244 1107 2245 1147
rect 2247 1107 2248 1147
rect 2252 1107 2253 1147
rect 2255 1107 2256 1147
rect 2304 1107 2305 1147
rect 2307 1107 2308 1147
rect 2312 1107 2313 1147
rect 2315 1107 2316 1147
rect 2364 1114 2365 1134
rect 2367 1114 2368 1134
rect 1023 1089 1083 1090
rect 1023 1086 1083 1087
rect 1023 1081 1083 1082
rect 1821 1084 1861 1085
rect 1023 1078 1083 1079
rect 1821 1081 1861 1082
rect 1821 1076 1861 1077
rect 1821 1073 1861 1074
rect 1212 1056 1272 1057
rect 1212 1053 1272 1054
rect 1212 1048 1272 1049
rect -539 937 -538 957
rect -536 937 -535 957
rect -487 951 -486 991
rect -484 951 -483 991
rect -479 951 -478 991
rect -476 951 -475 991
rect -427 951 -426 991
rect -424 951 -423 991
rect -419 951 -418 991
rect -416 951 -415 991
rect -367 958 -366 978
rect -364 958 -363 978
rect 1212 1045 1272 1046
rect 1212 1040 1272 1041
rect 288 1033 328 1034
rect 1212 1037 1272 1038
rect 288 1030 328 1031
rect 288 1025 328 1026
rect 288 1022 328 1023
rect 1029 1013 1069 1014
rect 1029 1010 1069 1011
rect 1029 1005 1069 1006
rect -208 947 -207 967
rect -205 947 -204 967
rect -156 961 -155 1001
rect -153 961 -152 1001
rect -148 961 -147 1001
rect -145 961 -144 1001
rect -96 961 -95 1001
rect -93 961 -92 1001
rect -88 961 -87 1001
rect -85 961 -84 1001
rect 1029 1002 1069 1003
rect 454 996 494 997
rect -36 968 -35 988
rect -33 968 -32 988
rect 454 993 494 994
rect 454 988 494 989
rect 454 985 494 986
rect 132 968 172 969
rect 1828 969 1868 970
rect 132 965 172 966
rect 132 960 172 961
rect 1828 966 1868 967
rect 1828 961 1868 962
rect 132 957 172 958
rect 1828 958 1868 959
rect 288 947 328 948
rect 288 944 328 945
rect 288 939 328 940
rect 288 936 328 937
rect 1015 931 1095 932
rect 1994 932 2034 933
rect 1015 928 1095 929
rect 1015 923 1095 924
rect 1994 929 2034 930
rect 1994 924 2034 925
rect 1015 920 1095 921
rect 1994 921 2034 922
rect 1015 915 1095 916
rect 1015 912 1095 913
rect 1015 907 1095 908
rect 1015 904 1095 905
rect 1672 904 1712 905
rect 1672 901 1712 902
rect 1672 896 1712 897
rect 1672 893 1712 894
rect 1234 882 1314 883
rect 1828 883 1868 884
rect 1234 879 1314 880
rect 1234 874 1314 875
rect 1828 880 1868 881
rect 1828 875 1868 876
rect 2185 873 2186 893
rect 2188 873 2189 893
rect 2237 887 2238 927
rect 2240 887 2241 927
rect 2245 887 2246 927
rect 2248 887 2249 927
rect 2297 887 2298 927
rect 2300 887 2301 927
rect 2305 887 2306 927
rect 2308 887 2309 927
rect 2357 894 2358 914
rect 2360 894 2361 914
rect 260 858 300 859
rect 260 855 300 856
rect 260 850 300 851
rect 260 847 300 848
rect 601 847 602 867
rect 604 847 605 867
rect 1234 871 1314 872
rect 1828 872 1868 873
rect 1234 866 1314 867
rect 1234 863 1314 864
rect 1234 858 1314 859
rect 1234 855 1314 856
rect 1019 834 1079 835
rect 1019 831 1079 832
rect 1019 826 1079 827
rect 1019 823 1079 824
rect 1019 818 1079 819
rect 1019 815 1079 816
rect 1025 761 1065 762
rect 1025 758 1065 759
rect 1025 753 1065 754
rect 1025 750 1065 751
rect -498 595 -497 615
rect -495 595 -494 615
rect -446 609 -445 649
rect -443 609 -442 649
rect -438 609 -437 649
rect -435 609 -434 649
rect -386 609 -385 649
rect -383 609 -382 649
rect -378 609 -377 649
rect -375 609 -374 649
rect -326 616 -325 636
rect -323 616 -322 636
rect 287 691 327 692
rect 287 688 327 689
rect 287 683 327 684
rect 287 680 327 681
rect -189 599 -188 619
rect -186 599 -185 619
rect -137 613 -136 653
rect -134 613 -133 653
rect -129 613 -128 653
rect -126 613 -125 653
rect -77 613 -76 653
rect -74 613 -73 653
rect -69 613 -68 653
rect -66 613 -65 653
rect 453 654 493 655
rect 453 651 493 652
rect 453 646 493 647
rect -17 620 -16 640
rect -14 620 -13 640
rect 453 643 493 644
rect 131 626 171 627
rect 131 623 171 624
rect 131 618 171 619
rect 131 615 171 616
rect 287 605 327 606
rect 287 602 327 603
rect 287 597 327 598
rect 287 594 327 595
rect 259 516 299 517
rect 259 513 299 514
rect 259 508 299 509
rect 259 505 299 506
rect 595 505 596 525
rect 598 505 599 525
rect 983 425 1063 426
rect 983 422 1063 423
rect 983 417 1063 418
rect 281 409 321 410
rect 281 406 321 407
rect 983 414 1063 415
rect 983 409 1063 410
rect 281 401 321 402
rect 281 398 321 399
rect 983 406 1063 407
rect 983 401 1063 402
rect 983 398 1063 399
rect 983 393 1063 394
rect 983 390 1063 391
rect 447 372 487 373
rect 447 369 487 370
rect 447 364 487 365
rect -579 264 -578 284
rect -576 264 -575 284
rect -527 278 -526 318
rect -524 278 -523 318
rect -519 278 -518 318
rect -516 278 -515 318
rect -467 278 -466 318
rect -464 278 -463 318
rect -459 278 -458 318
rect -456 278 -455 318
rect -407 285 -406 305
rect -404 285 -403 305
rect 447 361 487 362
rect 125 344 165 345
rect 125 341 165 342
rect 1267 340 1347 341
rect 125 336 165 337
rect 125 333 165 334
rect 1267 337 1347 338
rect 1267 332 1347 333
rect 281 323 321 324
rect 1267 329 1347 330
rect 1267 324 1347 325
rect -241 264 -240 284
rect -238 264 -237 284
rect -189 278 -188 318
rect -186 278 -185 318
rect -181 278 -180 318
rect -178 278 -177 318
rect -129 278 -128 318
rect -126 278 -125 318
rect -121 278 -120 318
rect -118 278 -117 318
rect 281 320 321 321
rect 281 315 321 316
rect 1267 321 1347 322
rect 1267 316 1347 317
rect 281 312 321 313
rect 1267 313 1347 314
rect 1267 308 1347 309
rect -69 285 -68 305
rect -66 285 -65 305
rect 1267 305 1347 306
rect 1005 264 1085 265
rect 1005 261 1085 262
rect 1005 256 1085 257
rect 1005 253 1085 254
rect 1005 248 1085 249
rect 1005 245 1085 246
rect 1005 240 1085 241
rect 253 234 293 235
rect 1005 237 1085 238
rect 253 231 293 232
rect 253 226 293 227
rect 253 223 293 224
rect 1628 212 1629 232
rect 1631 212 1632 232
rect 1680 226 1681 266
rect 1683 226 1684 266
rect 1688 226 1689 266
rect 1691 226 1692 266
rect 1740 226 1741 266
rect 1743 226 1744 266
rect 1748 226 1749 266
rect 1751 226 1752 266
rect 1800 233 1801 253
rect 1803 233 1804 253
rect 1012 120 1072 121
rect 1012 117 1072 118
rect 1012 112 1072 113
rect 1012 109 1072 110
rect 1012 104 1072 105
rect 1012 101 1072 102
rect 1029 30 1069 31
rect 1029 27 1069 28
rect 1029 22 1069 23
rect 1029 19 1069 20
<< pdiffusion >>
rect -120 1784 -119 1864
rect -117 1784 -116 1864
rect -112 1784 -111 1864
rect -109 1784 -108 1864
rect -68 1797 -67 1837
rect -65 1797 -64 1837
rect -8 1797 -7 1837
rect -5 1797 -4 1837
rect 52 1783 53 1823
rect 55 1783 56 1823
rect 682 1772 683 1852
rect 685 1772 686 1852
rect 690 1772 691 1852
rect 693 1772 694 1852
rect 734 1785 735 1825
rect 737 1785 738 1825
rect 794 1785 795 1825
rect 797 1785 798 1825
rect 854 1771 855 1811
rect 857 1771 858 1811
rect 256 1725 296 1726
rect 256 1722 296 1723
rect 256 1717 296 1718
rect 256 1714 296 1715
rect 422 1688 462 1689
rect 422 1685 462 1686
rect 422 1680 462 1681
rect 422 1677 462 1678
rect 100 1660 140 1661
rect 100 1657 140 1658
rect 100 1652 140 1653
rect 100 1649 140 1650
rect 256 1639 296 1640
rect 256 1636 296 1637
rect 256 1631 296 1632
rect 1764 1639 1804 1640
rect 1764 1636 1804 1637
rect 256 1628 296 1629
rect 1764 1631 1804 1632
rect 2180 1633 2181 1713
rect 2183 1633 2184 1713
rect 2188 1633 2189 1713
rect 2191 1633 2192 1713
rect 2232 1646 2233 1686
rect 2235 1646 2236 1686
rect 2292 1646 2293 1686
rect 2295 1646 2296 1686
rect 1764 1628 1804 1629
rect -190 1534 -189 1614
rect -187 1534 -186 1614
rect -182 1534 -181 1614
rect -179 1534 -178 1614
rect -138 1547 -137 1587
rect -135 1547 -134 1587
rect -78 1547 -77 1587
rect -75 1547 -74 1587
rect 619 1573 620 1613
rect 622 1573 623 1613
rect 1930 1602 1970 1603
rect 1930 1599 1970 1600
rect 1930 1594 1970 1595
rect 2352 1632 2353 1672
rect 2355 1632 2356 1672
rect 1930 1591 1970 1592
rect -18 1533 -17 1573
rect -15 1533 -14 1573
rect 1608 1574 1648 1575
rect 1608 1571 1648 1572
rect 1608 1566 1648 1567
rect 1608 1563 1648 1564
rect 228 1550 268 1551
rect 228 1547 268 1548
rect 228 1542 268 1543
rect 228 1539 268 1540
rect 1764 1553 1804 1554
rect 1764 1550 1804 1551
rect 1764 1545 1804 1546
rect 1764 1542 1804 1543
rect -515 1307 -514 1387
rect -512 1307 -511 1387
rect -507 1307 -506 1387
rect -504 1307 -503 1387
rect -463 1320 -462 1360
rect -460 1320 -459 1360
rect -403 1320 -402 1360
rect -400 1320 -399 1360
rect -343 1306 -342 1346
rect -340 1306 -339 1346
rect -158 1310 -157 1390
rect -155 1310 -154 1390
rect -150 1310 -149 1390
rect -147 1310 -146 1390
rect 263 1374 303 1375
rect 2184 1373 2185 1453
rect 2187 1373 2188 1453
rect 2192 1373 2193 1453
rect 2195 1373 2196 1453
rect 2236 1386 2237 1426
rect 2239 1386 2240 1426
rect 2296 1386 2297 1426
rect 2299 1386 2300 1426
rect 263 1371 303 1372
rect 263 1366 303 1367
rect 263 1363 303 1364
rect -106 1323 -105 1363
rect -103 1323 -102 1363
rect -46 1323 -45 1363
rect -43 1323 -42 1363
rect 1764 1364 1804 1365
rect 1764 1361 1804 1362
rect 1764 1356 1804 1357
rect 1764 1353 1804 1354
rect 14 1309 15 1349
rect 17 1309 18 1349
rect 429 1337 469 1338
rect 2356 1372 2357 1412
rect 2359 1372 2360 1412
rect 429 1334 469 1335
rect 429 1329 469 1330
rect 429 1326 469 1327
rect 1930 1327 1970 1328
rect 1930 1324 1970 1325
rect 1930 1319 1970 1320
rect 1930 1316 1970 1317
rect 107 1309 147 1310
rect 107 1306 147 1307
rect 107 1301 147 1302
rect 971 1304 1011 1305
rect 971 1301 1011 1302
rect 107 1298 147 1299
rect 971 1296 1011 1297
rect 1608 1299 1648 1300
rect 1608 1296 1648 1297
rect 971 1293 1011 1294
rect 263 1288 303 1289
rect 1608 1291 1648 1292
rect 1608 1288 1648 1289
rect 263 1285 303 1286
rect 263 1280 303 1281
rect 263 1277 303 1278
rect 1764 1278 1804 1279
rect 1764 1275 1804 1276
rect 1764 1270 1804 1271
rect 1764 1267 1804 1268
rect 622 1222 623 1262
rect 625 1222 626 1262
rect 1195 1239 1235 1240
rect 1195 1236 1235 1237
rect 1195 1231 1235 1232
rect 1195 1228 1235 1229
rect 235 1199 275 1200
rect 235 1196 275 1197
rect 235 1191 275 1192
rect 235 1188 275 1189
rect 1766 1170 1806 1171
rect 1766 1167 1806 1168
rect 1766 1162 1806 1163
rect 1766 1159 1806 1160
rect 2192 1149 2193 1229
rect 2195 1149 2196 1229
rect 2200 1149 2201 1229
rect 2203 1149 2204 1229
rect 2244 1162 2245 1202
rect 2247 1162 2248 1202
rect 2304 1162 2305 1202
rect 2307 1162 2308 1202
rect 1932 1133 1972 1134
rect 1932 1130 1972 1131
rect 1932 1125 1972 1126
rect 1932 1122 1972 1123
rect 2364 1148 2365 1188
rect 2367 1148 2368 1188
rect 1610 1105 1650 1106
rect 1610 1102 1650 1103
rect 965 1097 1005 1098
rect 965 1094 1005 1095
rect 965 1089 1005 1090
rect 1610 1097 1650 1098
rect 1610 1094 1650 1095
rect 965 1086 1005 1087
rect -539 993 -538 1073
rect -536 993 -535 1073
rect -531 993 -530 1073
rect -528 993 -527 1073
rect -487 1006 -486 1046
rect -484 1006 -483 1046
rect -427 1006 -426 1046
rect -424 1006 -423 1046
rect -367 992 -366 1032
rect -364 992 -363 1032
rect -208 1003 -207 1083
rect -205 1003 -204 1083
rect -200 1003 -199 1083
rect -197 1003 -196 1083
rect 965 1081 1005 1082
rect 1766 1084 1806 1085
rect 1766 1081 1806 1082
rect 965 1078 1005 1079
rect 1766 1076 1806 1077
rect 1766 1073 1806 1074
rect -156 1016 -155 1056
rect -153 1016 -152 1056
rect -96 1016 -95 1056
rect -93 1016 -92 1056
rect 1154 1056 1194 1057
rect 1154 1053 1194 1054
rect 1154 1048 1194 1049
rect 1154 1045 1194 1046
rect -36 1002 -35 1042
rect -33 1002 -32 1042
rect 233 1033 273 1034
rect 1154 1040 1194 1041
rect 1154 1037 1194 1038
rect 233 1030 273 1031
rect 233 1025 273 1026
rect 233 1022 273 1023
rect 974 1013 1014 1014
rect 974 1010 1014 1011
rect 974 1005 1014 1006
rect 974 1002 1014 1003
rect 399 996 439 997
rect 399 993 439 994
rect 399 988 439 989
rect 399 985 439 986
rect 77 968 117 969
rect 1773 969 1813 970
rect 1773 966 1813 967
rect 77 965 117 966
rect 77 960 117 961
rect 1773 961 1813 962
rect 1773 958 1813 959
rect 77 957 117 958
rect 233 947 273 948
rect 233 944 273 945
rect 233 939 273 940
rect 233 936 273 937
rect 951 931 991 932
rect 1939 932 1979 933
rect 1939 929 1979 930
rect 951 928 991 929
rect 601 881 602 921
rect 604 881 605 921
rect 951 923 991 924
rect 1939 924 1979 925
rect 2185 929 2186 1009
rect 2188 929 2189 1009
rect 2193 929 2194 1009
rect 2196 929 2197 1009
rect 2237 942 2238 982
rect 2240 942 2241 982
rect 2297 942 2298 982
rect 2300 942 2301 982
rect 1939 921 1979 922
rect 951 920 991 921
rect 951 915 991 916
rect 951 912 991 913
rect 951 907 991 908
rect 951 904 991 905
rect 1617 904 1657 905
rect 1617 901 1657 902
rect 1617 896 1657 897
rect 1617 893 1657 894
rect 2357 928 2358 968
rect 2360 928 2361 968
rect 1170 882 1210 883
rect 1773 883 1813 884
rect 1773 880 1813 881
rect 1170 879 1210 880
rect 1170 874 1210 875
rect 1773 875 1813 876
rect 1773 872 1813 873
rect 1170 871 1210 872
rect 205 858 245 859
rect 205 855 245 856
rect 205 850 245 851
rect 205 847 245 848
rect 1170 866 1210 867
rect 1170 863 1210 864
rect 1170 858 1210 859
rect 1170 855 1210 856
rect 961 834 1001 835
rect 961 831 1001 832
rect 961 826 1001 827
rect 961 823 1001 824
rect 961 818 1001 819
rect 961 815 1001 816
rect 970 761 1010 762
rect 970 758 1010 759
rect 970 753 1010 754
rect 970 750 1010 751
rect -498 651 -497 731
rect -495 651 -494 731
rect -490 651 -489 731
rect -487 651 -486 731
rect -446 664 -445 704
rect -443 664 -442 704
rect -386 664 -385 704
rect -383 664 -382 704
rect -326 650 -325 690
rect -323 650 -322 690
rect -189 655 -188 735
rect -186 655 -185 735
rect -181 655 -180 735
rect -178 655 -177 735
rect -137 668 -136 708
rect -134 668 -133 708
rect -77 668 -76 708
rect -74 668 -73 708
rect -17 654 -16 694
rect -14 654 -13 694
rect 232 691 272 692
rect 232 688 272 689
rect 232 683 272 684
rect 232 680 272 681
rect 398 654 438 655
rect 398 651 438 652
rect 398 646 438 647
rect 398 643 438 644
rect 76 626 116 627
rect 76 623 116 624
rect 76 618 116 619
rect 76 615 116 616
rect 232 605 272 606
rect 232 602 272 603
rect 232 597 272 598
rect 232 594 272 595
rect 595 539 596 579
rect 598 539 599 579
rect 204 516 244 517
rect 204 513 244 514
rect 204 508 244 509
rect 204 505 244 506
rect 919 425 959 426
rect 919 422 959 423
rect 919 417 959 418
rect 919 414 959 415
rect 226 409 266 410
rect 226 406 266 407
rect -579 320 -578 400
rect -576 320 -575 400
rect -571 320 -570 400
rect -568 320 -567 400
rect -527 333 -526 373
rect -524 333 -523 373
rect -467 333 -466 373
rect -464 333 -463 373
rect -407 319 -406 359
rect -404 319 -403 359
rect -241 320 -240 400
rect -238 320 -237 400
rect -233 320 -232 400
rect -230 320 -229 400
rect 226 401 266 402
rect 919 409 959 410
rect 919 406 959 407
rect 226 398 266 399
rect 919 401 959 402
rect 919 398 959 399
rect 919 393 959 394
rect 919 390 959 391
rect -189 333 -188 373
rect -186 333 -185 373
rect -129 333 -128 373
rect -126 333 -125 373
rect 392 372 432 373
rect 392 369 432 370
rect 392 364 432 365
rect 392 361 432 362
rect -69 319 -68 359
rect -66 319 -65 359
rect 70 344 110 345
rect 70 341 110 342
rect 70 336 110 337
rect 1203 340 1243 341
rect 1203 337 1243 338
rect 70 333 110 334
rect 1203 332 1243 333
rect 1203 329 1243 330
rect 226 323 266 324
rect 1203 324 1243 325
rect 1203 321 1243 322
rect 226 320 266 321
rect 226 315 266 316
rect 1203 316 1243 317
rect 1203 313 1243 314
rect 226 312 266 313
rect 1203 308 1243 309
rect 1203 305 1243 306
rect 941 264 981 265
rect 1628 268 1629 348
rect 1631 268 1632 348
rect 1636 268 1637 348
rect 1639 268 1640 348
rect 1680 281 1681 321
rect 1683 281 1684 321
rect 1740 281 1741 321
rect 1743 281 1744 321
rect 941 261 981 262
rect 941 256 981 257
rect 941 253 981 254
rect 941 248 981 249
rect 941 245 981 246
rect 198 234 238 235
rect 941 240 981 241
rect 941 237 981 238
rect 1800 267 1801 307
rect 1803 267 1804 307
rect 198 231 238 232
rect 198 226 238 227
rect 198 223 238 224
rect 954 120 994 121
rect 954 117 994 118
rect 954 112 994 113
rect 954 109 994 110
rect 954 104 994 105
rect 954 101 994 102
rect 974 30 1014 31
rect 974 27 1014 28
rect 974 22 1014 23
rect 974 19 1014 20
<< ndcontact >>
rect -124 1728 -120 1748
rect -116 1728 -112 1748
rect -72 1742 -68 1782
rect -64 1742 -60 1782
rect -56 1742 -52 1782
rect -12 1742 -8 1782
rect -4 1742 0 1782
rect 4 1742 8 1782
rect 48 1749 52 1769
rect 56 1749 60 1769
rect 311 1726 351 1730
rect 311 1718 351 1722
rect 678 1716 682 1736
rect 686 1716 690 1736
rect 730 1730 734 1770
rect 738 1730 742 1770
rect 746 1730 750 1770
rect 790 1730 794 1770
rect 798 1730 802 1770
rect 806 1730 810 1770
rect 850 1737 854 1757
rect 858 1737 862 1757
rect 311 1710 351 1714
rect 477 1689 517 1693
rect 477 1681 517 1685
rect 477 1673 517 1677
rect 155 1661 195 1665
rect 155 1653 195 1657
rect 155 1645 195 1649
rect 311 1640 351 1644
rect 1819 1640 1859 1644
rect 311 1632 351 1636
rect 1819 1632 1859 1636
rect 311 1624 351 1628
rect 1819 1624 1859 1628
rect 1985 1603 2025 1607
rect 1985 1595 2025 1599
rect 1985 1587 2025 1591
rect 1663 1575 1703 1579
rect 2176 1577 2180 1597
rect 2184 1577 2188 1597
rect 2228 1591 2232 1631
rect 2236 1591 2240 1631
rect 2244 1591 2248 1631
rect 2288 1591 2292 1631
rect 2296 1591 2300 1631
rect 2304 1591 2308 1631
rect 2348 1598 2352 1618
rect 2356 1598 2360 1618
rect 1663 1567 1703 1571
rect 1663 1559 1703 1563
rect 283 1551 323 1555
rect 283 1543 323 1547
rect 615 1539 619 1559
rect 623 1539 627 1559
rect 1819 1554 1859 1558
rect 1819 1546 1859 1550
rect 283 1535 323 1539
rect 1819 1538 1859 1542
rect -194 1478 -190 1498
rect -186 1478 -182 1498
rect -142 1492 -138 1532
rect -134 1492 -130 1532
rect -126 1492 -122 1532
rect -82 1492 -78 1532
rect -74 1492 -70 1532
rect -66 1492 -62 1532
rect -22 1499 -18 1519
rect -14 1499 -10 1519
rect 318 1375 358 1379
rect 318 1367 358 1371
rect 318 1359 358 1363
rect 1819 1365 1859 1369
rect 1819 1357 1859 1361
rect 1819 1349 1859 1353
rect -519 1251 -515 1271
rect -511 1251 -507 1271
rect -467 1265 -463 1305
rect -459 1265 -455 1305
rect -451 1265 -447 1305
rect -407 1265 -403 1305
rect -399 1265 -395 1305
rect -391 1265 -387 1305
rect -347 1272 -343 1292
rect -339 1272 -335 1292
rect 484 1338 524 1342
rect 484 1330 524 1334
rect 484 1322 524 1326
rect 1985 1328 2025 1332
rect 1985 1320 2025 1324
rect 2180 1317 2184 1337
rect 2188 1317 2192 1337
rect 2232 1331 2236 1371
rect 2240 1331 2244 1371
rect 2248 1331 2252 1371
rect 2292 1331 2296 1371
rect 2300 1331 2304 1371
rect 2308 1331 2312 1371
rect 2352 1338 2356 1358
rect 2360 1338 2364 1358
rect -162 1254 -158 1274
rect -154 1254 -150 1274
rect -110 1268 -106 1308
rect -102 1268 -98 1308
rect -94 1268 -90 1308
rect -50 1268 -46 1308
rect -42 1268 -38 1308
rect -34 1268 -30 1308
rect 162 1310 202 1314
rect 1985 1312 2025 1316
rect 162 1302 202 1306
rect 1026 1305 1066 1309
rect 10 1275 14 1295
rect 18 1275 22 1295
rect 162 1294 202 1298
rect 1026 1297 1066 1301
rect 1663 1300 1703 1304
rect 318 1289 358 1293
rect 1026 1289 1066 1293
rect 1663 1292 1703 1296
rect 318 1281 358 1285
rect 1663 1284 1703 1288
rect 318 1273 358 1277
rect 1819 1279 1859 1283
rect 1819 1271 1859 1275
rect 1819 1263 1859 1267
rect 1250 1240 1290 1244
rect 1250 1232 1290 1236
rect 1250 1224 1290 1228
rect 290 1200 330 1204
rect 290 1192 330 1196
rect 618 1188 622 1208
rect 626 1188 630 1208
rect 290 1184 330 1188
rect 1821 1171 1861 1175
rect 1821 1163 1861 1167
rect 1821 1155 1861 1159
rect 1987 1134 2027 1138
rect 1987 1126 2027 1130
rect 1987 1118 2027 1122
rect 1665 1106 1705 1110
rect 1023 1098 1083 1102
rect 1665 1098 1705 1102
rect 1023 1090 1083 1094
rect 1665 1090 1705 1094
rect 2188 1093 2192 1113
rect 2196 1093 2200 1113
rect 2240 1107 2244 1147
rect 2248 1107 2252 1147
rect 2256 1107 2260 1147
rect 2300 1107 2304 1147
rect 2308 1107 2312 1147
rect 2316 1107 2320 1147
rect 2360 1114 2364 1134
rect 2368 1114 2372 1134
rect 1023 1082 1083 1086
rect 1821 1085 1861 1089
rect 1023 1074 1083 1078
rect 1821 1077 1861 1081
rect 1821 1069 1861 1073
rect 1212 1057 1272 1061
rect 1212 1049 1272 1053
rect -543 937 -539 957
rect -535 937 -531 957
rect -491 951 -487 991
rect -483 951 -479 991
rect -475 951 -471 991
rect -431 951 -427 991
rect -423 951 -419 991
rect -415 951 -411 991
rect -371 958 -367 978
rect -363 958 -359 978
rect 288 1034 328 1038
rect 1212 1041 1272 1045
rect 1212 1033 1272 1037
rect 288 1026 328 1030
rect 288 1018 328 1022
rect 1029 1014 1069 1018
rect 1029 1006 1069 1010
rect -212 947 -208 967
rect -204 947 -200 967
rect -160 961 -156 1001
rect -152 961 -148 1001
rect -144 961 -140 1001
rect -100 961 -96 1001
rect -92 961 -88 1001
rect -84 961 -80 1001
rect 454 997 494 1001
rect 1029 998 1069 1002
rect -40 968 -36 988
rect -32 968 -28 988
rect 454 989 494 993
rect 454 981 494 985
rect 132 969 172 973
rect 1828 970 1868 974
rect 132 961 172 965
rect 1828 962 1868 966
rect 132 953 172 957
rect 1828 954 1868 958
rect 288 948 328 952
rect 288 940 328 944
rect 288 932 328 936
rect 1015 932 1095 936
rect 1994 933 2034 937
rect 1015 924 1095 928
rect 1994 925 2034 929
rect 1015 916 1095 920
rect 1994 917 2034 921
rect 1015 908 1095 912
rect 1015 900 1095 904
rect 1672 905 1712 909
rect 1672 897 1712 901
rect 1672 889 1712 893
rect 1234 883 1314 887
rect 1828 884 1868 888
rect 1234 875 1314 879
rect 1828 876 1868 880
rect 2181 873 2185 893
rect 2189 873 2193 893
rect 2233 887 2237 927
rect 2241 887 2245 927
rect 2249 887 2253 927
rect 2293 887 2297 927
rect 2301 887 2305 927
rect 2309 887 2313 927
rect 2353 894 2357 914
rect 2361 894 2365 914
rect 260 859 300 863
rect 260 851 300 855
rect 597 847 601 867
rect 605 847 609 867
rect 1234 867 1314 871
rect 1828 868 1868 872
rect 1234 859 1314 863
rect 1234 851 1314 855
rect 260 843 300 847
rect 1019 835 1079 839
rect 1019 827 1079 831
rect 1019 819 1079 823
rect 1019 811 1079 815
rect 1025 762 1065 766
rect 1025 754 1065 758
rect 1025 746 1065 750
rect -502 595 -498 615
rect -494 595 -490 615
rect -450 609 -446 649
rect -442 609 -438 649
rect -434 609 -430 649
rect -390 609 -386 649
rect -382 609 -378 649
rect -374 609 -370 649
rect -330 616 -326 636
rect -322 616 -318 636
rect 287 692 327 696
rect 287 684 327 688
rect 287 676 327 680
rect -193 599 -189 619
rect -185 599 -181 619
rect -141 613 -137 653
rect -133 613 -129 653
rect -125 613 -121 653
rect -81 613 -77 653
rect -73 613 -69 653
rect -65 613 -61 653
rect 453 655 493 659
rect 453 647 493 651
rect -21 620 -17 640
rect -13 620 -9 640
rect 453 639 493 643
rect 131 627 171 631
rect 131 619 171 623
rect 131 611 171 615
rect 287 606 327 610
rect 287 598 327 602
rect 287 590 327 594
rect 259 517 299 521
rect 259 509 299 513
rect 591 505 595 525
rect 599 505 603 525
rect 259 501 299 505
rect 983 426 1063 430
rect 983 418 1063 422
rect 281 410 321 414
rect 983 410 1063 414
rect 281 402 321 406
rect 983 402 1063 406
rect 281 394 321 398
rect 983 394 1063 398
rect 983 386 1063 390
rect 447 373 487 377
rect 447 365 487 369
rect -583 264 -579 284
rect -575 264 -571 284
rect -531 278 -527 318
rect -523 278 -519 318
rect -515 278 -511 318
rect -471 278 -467 318
rect -463 278 -459 318
rect -455 278 -451 318
rect -411 285 -407 305
rect -403 285 -399 305
rect 447 357 487 361
rect 125 345 165 349
rect 125 337 165 341
rect 1267 341 1347 345
rect 125 329 165 333
rect 1267 333 1347 337
rect 281 324 321 328
rect 1267 325 1347 329
rect -245 264 -241 284
rect -237 264 -233 284
rect -193 278 -189 318
rect -185 278 -181 318
rect -177 278 -173 318
rect -133 278 -129 318
rect -125 278 -121 318
rect -117 278 -113 318
rect 281 316 321 320
rect 1267 317 1347 321
rect 281 308 321 312
rect 1267 309 1347 313
rect -73 285 -69 305
rect -65 285 -61 305
rect 1267 301 1347 305
rect 1005 265 1085 269
rect 1005 257 1085 261
rect 1005 249 1085 253
rect 253 235 293 239
rect 1005 241 1085 245
rect 1005 233 1085 237
rect 253 227 293 231
rect 253 219 293 223
rect 1624 212 1628 232
rect 1632 212 1636 232
rect 1676 226 1680 266
rect 1684 226 1688 266
rect 1692 226 1696 266
rect 1736 226 1740 266
rect 1744 226 1748 266
rect 1752 226 1756 266
rect 1796 233 1800 253
rect 1804 233 1808 253
rect 1012 121 1072 125
rect 1012 113 1072 117
rect 1012 105 1072 109
rect 1012 97 1072 101
rect 1029 31 1069 35
rect 1029 23 1069 27
rect 1029 15 1069 19
<< pdcontact >>
rect -124 1784 -120 1864
rect -116 1784 -112 1864
rect -108 1784 -104 1864
rect -72 1797 -68 1837
rect -64 1797 -60 1837
rect -12 1797 -8 1837
rect -4 1797 0 1837
rect 48 1783 52 1823
rect 56 1783 60 1823
rect 678 1772 682 1852
rect 686 1772 690 1852
rect 694 1772 698 1852
rect 730 1785 734 1825
rect 738 1785 742 1825
rect 790 1785 794 1825
rect 798 1785 802 1825
rect 850 1771 854 1811
rect 858 1771 862 1811
rect 256 1726 296 1730
rect 256 1718 296 1722
rect 256 1710 296 1714
rect 422 1689 462 1693
rect 422 1681 462 1685
rect 422 1673 462 1677
rect 100 1661 140 1665
rect 100 1653 140 1657
rect 100 1645 140 1649
rect 256 1640 296 1644
rect 1764 1640 1804 1644
rect 256 1632 296 1636
rect 1764 1632 1804 1636
rect 256 1624 296 1628
rect 2176 1633 2180 1713
rect 2184 1633 2188 1713
rect 2192 1633 2196 1713
rect 2228 1646 2232 1686
rect 2236 1646 2240 1686
rect 2288 1646 2292 1686
rect 2296 1646 2300 1686
rect 1764 1624 1804 1628
rect -194 1534 -190 1614
rect -186 1534 -182 1614
rect -178 1534 -174 1614
rect -142 1547 -138 1587
rect -134 1547 -130 1587
rect -82 1547 -78 1587
rect -74 1547 -70 1587
rect 615 1573 619 1613
rect 623 1573 627 1613
rect 1930 1603 1970 1607
rect 1930 1595 1970 1599
rect 2348 1632 2352 1672
rect 2356 1632 2360 1672
rect 1930 1587 1970 1591
rect 1608 1575 1648 1579
rect -22 1533 -18 1573
rect -14 1533 -10 1573
rect 1608 1567 1648 1571
rect 1608 1559 1648 1563
rect 228 1551 268 1555
rect 228 1543 268 1547
rect 228 1535 268 1539
rect 1764 1554 1804 1558
rect 1764 1546 1804 1550
rect 1764 1538 1804 1542
rect -519 1307 -515 1387
rect -511 1307 -507 1387
rect -503 1307 -499 1387
rect -467 1320 -463 1360
rect -459 1320 -455 1360
rect -407 1320 -403 1360
rect -399 1320 -395 1360
rect -347 1306 -343 1346
rect -339 1306 -335 1346
rect -162 1310 -158 1390
rect -154 1310 -150 1390
rect -146 1310 -142 1390
rect 263 1375 303 1379
rect 2180 1373 2184 1453
rect 2188 1373 2192 1453
rect 2196 1373 2200 1453
rect 2232 1386 2236 1426
rect 2240 1386 2244 1426
rect 2292 1386 2296 1426
rect 2300 1386 2304 1426
rect 263 1367 303 1371
rect 1764 1365 1804 1369
rect -110 1323 -106 1363
rect -102 1323 -98 1363
rect -50 1323 -46 1363
rect -42 1323 -38 1363
rect 263 1359 303 1363
rect 1764 1357 1804 1361
rect 1764 1349 1804 1353
rect 10 1309 14 1349
rect 18 1309 22 1349
rect 429 1338 469 1342
rect 2352 1372 2356 1412
rect 2360 1372 2364 1412
rect 429 1330 469 1334
rect 1930 1328 1970 1332
rect 429 1322 469 1326
rect 1930 1320 1970 1324
rect 107 1310 147 1314
rect 1930 1312 1970 1316
rect 107 1302 147 1306
rect 971 1305 1011 1309
rect 107 1294 147 1298
rect 971 1297 1011 1301
rect 1608 1300 1648 1304
rect 263 1289 303 1293
rect 971 1289 1011 1293
rect 1608 1292 1648 1296
rect 263 1281 303 1285
rect 1608 1284 1648 1288
rect 1764 1279 1804 1283
rect 263 1273 303 1277
rect 1764 1271 1804 1275
rect 1764 1263 1804 1267
rect 618 1222 622 1262
rect 626 1222 630 1262
rect 1195 1240 1235 1244
rect 1195 1232 1235 1236
rect 1195 1224 1235 1228
rect 235 1200 275 1204
rect 235 1192 275 1196
rect 235 1184 275 1188
rect 1766 1171 1806 1175
rect 1766 1163 1806 1167
rect 1766 1155 1806 1159
rect 2188 1149 2192 1229
rect 2196 1149 2200 1229
rect 2204 1149 2208 1229
rect 2240 1162 2244 1202
rect 2248 1162 2252 1202
rect 2300 1162 2304 1202
rect 2308 1162 2312 1202
rect 1932 1134 1972 1138
rect 1932 1126 1972 1130
rect 1932 1118 1972 1122
rect 2360 1148 2364 1188
rect 2368 1148 2372 1188
rect 1610 1106 1650 1110
rect 965 1098 1005 1102
rect 1610 1098 1650 1102
rect 965 1090 1005 1094
rect 1610 1090 1650 1094
rect -543 993 -539 1073
rect -535 993 -531 1073
rect -527 993 -523 1073
rect -491 1006 -487 1046
rect -483 1006 -479 1046
rect -431 1006 -427 1046
rect -423 1006 -419 1046
rect -371 992 -367 1032
rect -363 992 -359 1032
rect -212 1003 -208 1083
rect -204 1003 -200 1083
rect -196 1003 -192 1083
rect 965 1082 1005 1086
rect 1766 1085 1806 1089
rect 965 1074 1005 1078
rect 1766 1077 1806 1081
rect 1766 1069 1806 1073
rect 1154 1057 1194 1061
rect -160 1016 -156 1056
rect -152 1016 -148 1056
rect -100 1016 -96 1056
rect -92 1016 -88 1056
rect 1154 1049 1194 1053
rect -40 1002 -36 1042
rect -32 1002 -28 1042
rect 1154 1041 1194 1045
rect 233 1034 273 1038
rect 1154 1033 1194 1037
rect 233 1026 273 1030
rect 233 1018 273 1022
rect 974 1014 1014 1018
rect 974 1006 1014 1010
rect 399 997 439 1001
rect 974 998 1014 1002
rect 399 989 439 993
rect 399 981 439 985
rect 77 969 117 973
rect 1773 970 1813 974
rect 77 961 117 965
rect 1773 962 1813 966
rect 77 953 117 957
rect 1773 954 1813 958
rect 233 948 273 952
rect 233 940 273 944
rect 233 932 273 936
rect 951 932 991 936
rect 1939 933 1979 937
rect 951 924 991 928
rect 597 881 601 921
rect 605 881 609 921
rect 1939 925 1979 929
rect 2181 929 2185 1009
rect 2189 929 2193 1009
rect 2197 929 2201 1009
rect 2233 942 2237 982
rect 2241 942 2245 982
rect 2293 942 2297 982
rect 2301 942 2305 982
rect 951 916 991 920
rect 1939 917 1979 921
rect 951 908 991 912
rect 1617 905 1657 909
rect 951 900 991 904
rect 1617 897 1657 901
rect 1617 889 1657 893
rect 2353 928 2357 968
rect 2361 928 2365 968
rect 1170 883 1210 887
rect 1773 884 1813 888
rect 1170 875 1210 879
rect 1773 876 1813 880
rect 1170 867 1210 871
rect 205 859 245 863
rect 205 851 245 855
rect 205 843 245 847
rect 1773 868 1813 872
rect 1170 859 1210 863
rect 1170 851 1210 855
rect 961 835 1001 839
rect 961 827 1001 831
rect 961 819 1001 823
rect 961 811 1001 815
rect 970 762 1010 766
rect 970 754 1010 758
rect 970 746 1010 750
rect -502 651 -498 731
rect -494 651 -490 731
rect -486 651 -482 731
rect -450 664 -446 704
rect -442 664 -438 704
rect -390 664 -386 704
rect -382 664 -378 704
rect -330 650 -326 690
rect -322 650 -318 690
rect -193 655 -189 735
rect -185 655 -181 735
rect -177 655 -173 735
rect -141 668 -137 708
rect -133 668 -129 708
rect -81 668 -77 708
rect -73 668 -69 708
rect -21 654 -17 694
rect -13 654 -9 694
rect 232 692 272 696
rect 232 684 272 688
rect 232 676 272 680
rect 398 655 438 659
rect 398 647 438 651
rect 398 639 438 643
rect 76 627 116 631
rect 76 619 116 623
rect 76 611 116 615
rect 232 606 272 610
rect 232 598 272 602
rect 232 590 272 594
rect 591 539 595 579
rect 599 539 603 579
rect 204 517 244 521
rect 204 509 244 513
rect 204 501 244 505
rect 919 426 959 430
rect 919 418 959 422
rect 226 410 266 414
rect 919 410 959 414
rect 226 402 266 406
rect -583 320 -579 400
rect -575 320 -571 400
rect -567 320 -563 400
rect -531 333 -527 373
rect -523 333 -519 373
rect -471 333 -467 373
rect -463 333 -459 373
rect -411 319 -407 359
rect -403 319 -399 359
rect -245 320 -241 400
rect -237 320 -233 400
rect -229 320 -225 400
rect 919 402 959 406
rect 226 394 266 398
rect 919 394 959 398
rect 919 386 959 390
rect 392 373 432 377
rect -193 333 -189 373
rect -185 333 -181 373
rect -133 333 -129 373
rect -125 333 -121 373
rect 392 365 432 369
rect -73 319 -69 359
rect -65 319 -61 359
rect 392 357 432 361
rect 70 345 110 349
rect 70 337 110 341
rect 1203 341 1243 345
rect 70 329 110 333
rect 1203 333 1243 337
rect 226 324 266 328
rect 1203 325 1243 329
rect 226 316 266 320
rect 1203 317 1243 321
rect 226 308 266 312
rect 1203 309 1243 313
rect 1203 301 1243 305
rect 941 265 981 269
rect 1624 268 1628 348
rect 1632 268 1636 348
rect 1640 268 1644 348
rect 1676 281 1680 321
rect 1684 281 1688 321
rect 1736 281 1740 321
rect 1744 281 1748 321
rect 941 257 981 261
rect 941 249 981 253
rect 941 241 981 245
rect 198 235 238 239
rect 941 233 981 237
rect 1796 267 1800 307
rect 1804 267 1808 307
rect 198 227 238 231
rect 198 219 238 223
rect 954 121 994 125
rect 954 113 994 117
rect 954 105 994 109
rect 954 97 994 101
rect 974 31 1014 35
rect 974 23 1014 27
rect 974 15 1014 19
<< polysilicon >>
rect -119 1864 -117 1877
rect -111 1864 -109 1877
rect 683 1852 685 1865
rect 691 1852 693 1865
rect -67 1837 -65 1848
rect -7 1837 -5 1848
rect 53 1823 55 1826
rect -119 1748 -117 1784
rect -111 1773 -109 1784
rect -67 1782 -65 1797
rect -59 1782 -57 1785
rect -7 1782 -5 1797
rect 1 1782 3 1785
rect 53 1769 55 1783
rect 735 1825 737 1836
rect 795 1825 797 1836
rect 855 1811 857 1814
rect 53 1746 55 1749
rect -67 1738 -65 1742
rect -59 1738 -57 1742
rect -7 1738 -5 1742
rect 1 1738 3 1742
rect 683 1736 685 1772
rect 691 1761 693 1772
rect 735 1770 737 1785
rect 743 1770 745 1773
rect 795 1770 797 1785
rect 803 1770 805 1773
rect -119 1724 -117 1728
rect 245 1723 256 1725
rect 296 1723 311 1725
rect 351 1723 355 1725
rect 245 1715 256 1717
rect 296 1715 311 1717
rect 351 1715 355 1717
rect 855 1757 857 1771
rect 855 1734 857 1737
rect 735 1726 737 1730
rect 743 1726 745 1730
rect 795 1726 797 1730
rect 803 1726 805 1730
rect 683 1712 685 1716
rect 2181 1713 2183 1726
rect 2189 1713 2191 1726
rect 411 1686 422 1688
rect 462 1686 477 1688
rect 517 1686 521 1688
rect 411 1678 422 1680
rect 462 1678 477 1680
rect 517 1678 521 1680
rect 89 1658 100 1660
rect 140 1658 155 1660
rect 195 1658 199 1660
rect 89 1650 100 1652
rect 140 1650 155 1652
rect 195 1650 199 1652
rect 245 1637 256 1639
rect 296 1637 311 1639
rect 351 1637 355 1639
rect 1753 1637 1764 1639
rect 1804 1637 1819 1639
rect 1859 1637 1863 1639
rect 245 1629 256 1631
rect 296 1629 311 1631
rect 351 1629 355 1631
rect -189 1614 -187 1627
rect -181 1614 -179 1627
rect 2233 1686 2235 1697
rect 2293 1686 2295 1697
rect 2353 1672 2355 1675
rect 1753 1629 1764 1631
rect 1804 1629 1819 1631
rect 1859 1629 1863 1631
rect 620 1613 622 1616
rect -137 1587 -135 1598
rect -77 1587 -75 1598
rect -17 1573 -15 1576
rect 1919 1600 1930 1602
rect 1970 1600 1985 1602
rect 2025 1600 2029 1602
rect 2181 1597 2183 1633
rect 2189 1622 2191 1633
rect 2233 1631 2235 1646
rect 2241 1631 2243 1634
rect 2293 1631 2295 1646
rect 2301 1631 2303 1634
rect 1919 1592 1930 1594
rect 1970 1592 1985 1594
rect 2025 1592 2029 1594
rect -189 1498 -187 1534
rect -181 1523 -179 1534
rect -137 1532 -135 1547
rect -129 1532 -127 1535
rect -77 1532 -75 1547
rect -69 1532 -67 1535
rect 620 1559 622 1573
rect 2353 1618 2355 1632
rect 2353 1595 2355 1598
rect 2233 1587 2235 1591
rect 2241 1587 2243 1591
rect 2293 1587 2295 1591
rect 2301 1587 2303 1591
rect 1597 1572 1608 1574
rect 1648 1572 1663 1574
rect 1703 1572 1707 1574
rect 2181 1573 2183 1577
rect 1597 1564 1608 1566
rect 1648 1564 1663 1566
rect 1703 1564 1707 1566
rect 217 1548 228 1550
rect 268 1548 283 1550
rect 323 1548 327 1550
rect 217 1540 228 1542
rect 268 1540 283 1542
rect 323 1540 327 1542
rect 1753 1551 1764 1553
rect 1804 1551 1819 1553
rect 1859 1551 1863 1553
rect 1753 1543 1764 1545
rect 1804 1543 1819 1545
rect 1859 1543 1863 1545
rect 620 1536 622 1539
rect -17 1519 -15 1533
rect -17 1496 -15 1499
rect -137 1488 -135 1492
rect -129 1488 -127 1492
rect -77 1488 -75 1492
rect -69 1488 -67 1492
rect -189 1474 -187 1478
rect 2185 1453 2187 1466
rect 2193 1453 2195 1466
rect -514 1387 -512 1400
rect -506 1387 -504 1400
rect -157 1390 -155 1403
rect -149 1390 -147 1403
rect -462 1360 -460 1371
rect -402 1360 -400 1371
rect -342 1346 -340 1349
rect -514 1271 -512 1307
rect -506 1296 -504 1307
rect -462 1305 -460 1320
rect -454 1305 -452 1308
rect -402 1305 -400 1320
rect -394 1305 -392 1308
rect -105 1363 -103 1374
rect -45 1363 -43 1374
rect 252 1372 263 1374
rect 303 1372 318 1374
rect 358 1372 362 1374
rect 2237 1426 2239 1437
rect 2297 1426 2299 1437
rect 2357 1412 2359 1415
rect 252 1364 263 1366
rect 303 1364 318 1366
rect 358 1364 362 1366
rect 1753 1362 1764 1364
rect 1804 1362 1819 1364
rect 1859 1362 1863 1364
rect 1753 1354 1764 1356
rect 1804 1354 1819 1356
rect 1859 1354 1863 1356
rect 15 1349 17 1352
rect -342 1292 -340 1306
rect -157 1274 -155 1310
rect -149 1299 -147 1310
rect -105 1308 -103 1323
rect -97 1308 -95 1311
rect -45 1308 -43 1323
rect -37 1308 -35 1311
rect 2185 1337 2187 1373
rect 2193 1362 2195 1373
rect 2237 1371 2239 1386
rect 2245 1371 2247 1374
rect 2297 1371 2299 1386
rect 2305 1371 2307 1374
rect 418 1335 429 1337
rect 469 1335 484 1337
rect 524 1335 528 1337
rect 418 1327 429 1329
rect 469 1327 484 1329
rect 524 1327 528 1329
rect 1919 1325 1930 1327
rect 1970 1325 1985 1327
rect 2025 1325 2029 1327
rect 1919 1317 1930 1319
rect 1970 1317 1985 1319
rect 2025 1317 2029 1319
rect 2357 1358 2359 1372
rect 2357 1335 2359 1338
rect 2237 1327 2239 1331
rect 2245 1327 2247 1331
rect 2297 1327 2299 1331
rect 2305 1327 2307 1331
rect -342 1269 -340 1272
rect -462 1261 -460 1265
rect -454 1261 -452 1265
rect -402 1261 -400 1265
rect -394 1261 -392 1265
rect 15 1295 17 1309
rect 2185 1313 2187 1317
rect 96 1307 107 1309
rect 147 1307 162 1309
rect 202 1307 206 1309
rect 960 1302 971 1304
rect 1011 1302 1026 1304
rect 1066 1302 1070 1304
rect 96 1299 107 1301
rect 147 1299 162 1301
rect 202 1299 206 1301
rect 1597 1297 1608 1299
rect 1648 1297 1663 1299
rect 1703 1297 1707 1299
rect 960 1294 971 1296
rect 1011 1294 1026 1296
rect 1066 1294 1070 1296
rect 1597 1289 1608 1291
rect 1648 1289 1663 1291
rect 1703 1289 1707 1291
rect 252 1286 263 1288
rect 303 1286 318 1288
rect 358 1286 362 1288
rect 252 1278 263 1280
rect 303 1278 318 1280
rect 358 1278 362 1280
rect 15 1272 17 1275
rect 1753 1276 1764 1278
rect 1804 1276 1819 1278
rect 1859 1276 1863 1278
rect -105 1264 -103 1268
rect -97 1264 -95 1268
rect -45 1264 -43 1268
rect -37 1264 -35 1268
rect 1753 1268 1764 1270
rect 1804 1268 1819 1270
rect 1859 1268 1863 1270
rect 623 1262 625 1265
rect -514 1247 -512 1251
rect -157 1250 -155 1254
rect 1184 1237 1195 1239
rect 1235 1237 1250 1239
rect 1290 1237 1294 1239
rect 1184 1229 1195 1231
rect 1235 1229 1250 1231
rect 1290 1229 1294 1231
rect 2193 1229 2195 1242
rect 2201 1229 2203 1242
rect 623 1208 625 1222
rect 224 1197 235 1199
rect 275 1197 290 1199
rect 330 1197 334 1199
rect 224 1189 235 1191
rect 275 1189 290 1191
rect 330 1189 334 1191
rect 623 1185 625 1188
rect 1755 1168 1766 1170
rect 1806 1168 1821 1170
rect 1861 1168 1865 1170
rect 1755 1160 1766 1162
rect 1806 1160 1821 1162
rect 1861 1160 1865 1162
rect 2245 1202 2247 1213
rect 2305 1202 2307 1213
rect 2365 1188 2367 1191
rect 1921 1131 1932 1133
rect 1972 1131 1987 1133
rect 2027 1131 2031 1133
rect 1921 1123 1932 1125
rect 1972 1123 1987 1125
rect 2027 1123 2031 1125
rect 2193 1113 2195 1149
rect 2201 1138 2203 1149
rect 2245 1147 2247 1162
rect 2253 1147 2255 1150
rect 2305 1147 2307 1162
rect 2313 1147 2315 1150
rect 1599 1103 1610 1105
rect 1650 1103 1665 1105
rect 1705 1103 1709 1105
rect -538 1073 -536 1086
rect -530 1073 -528 1086
rect -207 1083 -205 1096
rect -199 1083 -197 1096
rect 954 1095 965 1097
rect 1005 1095 1023 1097
rect 1083 1095 1088 1097
rect 1599 1095 1610 1097
rect 1650 1095 1665 1097
rect 1705 1095 1709 1097
rect 2365 1134 2367 1148
rect 2365 1111 2367 1114
rect 2245 1103 2247 1107
rect 2253 1103 2255 1107
rect 2305 1103 2307 1107
rect 2313 1103 2315 1107
rect 2193 1089 2195 1093
rect 954 1087 965 1089
rect 1005 1087 1023 1089
rect 1083 1087 1088 1089
rect -486 1046 -484 1057
rect -426 1046 -424 1057
rect -366 1032 -364 1035
rect -538 957 -536 993
rect -530 982 -528 993
rect -486 991 -484 1006
rect -478 991 -476 994
rect -426 991 -424 1006
rect -418 991 -416 994
rect 1755 1082 1766 1084
rect 1806 1082 1821 1084
rect 1861 1082 1865 1084
rect 954 1079 965 1081
rect 1005 1079 1023 1081
rect 1083 1079 1088 1081
rect 1755 1074 1766 1076
rect 1806 1074 1821 1076
rect 1861 1074 1865 1076
rect -155 1056 -153 1067
rect -95 1056 -93 1067
rect 1143 1054 1154 1056
rect 1194 1054 1212 1056
rect 1272 1054 1277 1056
rect 1143 1046 1154 1048
rect 1194 1046 1212 1048
rect 1272 1046 1277 1048
rect -35 1042 -33 1045
rect -366 978 -364 992
rect -207 967 -205 1003
rect -199 992 -197 1003
rect -155 1001 -153 1016
rect -147 1001 -145 1004
rect -95 1001 -93 1016
rect -87 1001 -85 1004
rect 1143 1038 1154 1040
rect 1194 1038 1212 1040
rect 1272 1038 1277 1040
rect 222 1031 233 1033
rect 273 1031 288 1033
rect 328 1031 332 1033
rect 222 1023 233 1025
rect 273 1023 288 1025
rect 328 1023 332 1025
rect 963 1011 974 1013
rect 1014 1011 1029 1013
rect 1069 1011 1073 1013
rect 2186 1009 2188 1022
rect 2194 1009 2196 1022
rect 963 1003 974 1005
rect 1014 1003 1029 1005
rect 1069 1003 1073 1005
rect -366 955 -364 958
rect -486 947 -484 951
rect -478 947 -476 951
rect -426 947 -424 951
rect -418 947 -416 951
rect -35 988 -33 1002
rect 388 994 399 996
rect 439 994 454 996
rect 494 994 498 996
rect 388 986 399 988
rect 439 986 454 988
rect 494 986 498 988
rect -35 965 -33 968
rect 66 966 77 968
rect 117 966 132 968
rect 172 966 176 968
rect 1762 967 1773 969
rect 1813 967 1828 969
rect 1868 967 1872 969
rect -155 957 -153 961
rect -147 957 -145 961
rect -95 957 -93 961
rect -87 957 -85 961
rect 66 958 77 960
rect 117 958 132 960
rect 172 958 176 960
rect 1762 959 1773 961
rect 1813 959 1828 961
rect 1868 959 1872 961
rect -207 943 -205 947
rect 222 945 233 947
rect 273 945 288 947
rect 328 945 332 947
rect -538 933 -536 937
rect 222 937 233 939
rect 273 937 288 939
rect 328 937 332 939
rect 940 929 951 931
rect 991 929 1015 931
rect 1095 929 1098 931
rect 1928 930 1939 932
rect 1979 930 1994 932
rect 2034 930 2038 932
rect 602 921 604 924
rect 940 921 951 923
rect 991 921 1015 923
rect 1095 921 1098 923
rect 2238 982 2240 993
rect 2298 982 2300 993
rect 2358 968 2360 971
rect 1928 922 1939 924
rect 1979 922 1994 924
rect 2034 922 2038 924
rect 940 913 951 915
rect 991 913 1015 915
rect 1095 913 1098 915
rect 940 905 951 907
rect 991 905 1015 907
rect 1095 905 1098 907
rect 1606 902 1617 904
rect 1657 902 1672 904
rect 1712 902 1716 904
rect 1606 894 1617 896
rect 1657 894 1672 896
rect 1712 894 1716 896
rect 2186 893 2188 929
rect 2194 918 2196 929
rect 2238 927 2240 942
rect 2246 927 2248 930
rect 2298 927 2300 942
rect 2306 927 2308 930
rect 602 867 604 881
rect 1159 880 1170 882
rect 1210 880 1234 882
rect 1314 880 1317 882
rect 1762 881 1773 883
rect 1813 881 1828 883
rect 1868 881 1872 883
rect 1159 872 1170 874
rect 1210 872 1234 874
rect 1314 872 1317 874
rect 1762 873 1773 875
rect 1813 873 1828 875
rect 1868 873 1872 875
rect 2358 914 2360 928
rect 2358 891 2360 894
rect 2238 883 2240 887
rect 2246 883 2248 887
rect 2298 883 2300 887
rect 2306 883 2308 887
rect 194 856 205 858
rect 245 856 260 858
rect 300 856 304 858
rect 194 848 205 850
rect 245 848 260 850
rect 300 848 304 850
rect 2186 869 2188 873
rect 1159 864 1170 866
rect 1210 864 1234 866
rect 1314 864 1317 866
rect 1159 856 1170 858
rect 1210 856 1234 858
rect 1314 856 1317 858
rect 602 844 604 847
rect 950 832 961 834
rect 1001 832 1019 834
rect 1079 832 1084 834
rect 950 824 961 826
rect 1001 824 1019 826
rect 1079 824 1084 826
rect 950 816 961 818
rect 1001 816 1019 818
rect 1079 816 1084 818
rect 959 759 970 761
rect 1010 759 1025 761
rect 1065 759 1069 761
rect 959 751 970 753
rect 1010 751 1025 753
rect 1065 751 1069 753
rect -497 731 -495 744
rect -489 731 -487 744
rect -188 735 -186 748
rect -180 735 -178 748
rect -445 704 -443 715
rect -385 704 -383 715
rect -325 690 -323 693
rect -497 615 -495 651
rect -489 640 -487 651
rect -445 649 -443 664
rect -437 649 -435 652
rect -385 649 -383 664
rect -377 649 -375 652
rect -136 708 -134 719
rect -76 708 -74 719
rect -16 694 -14 697
rect -325 636 -323 650
rect -188 619 -186 655
rect -180 644 -178 655
rect -136 653 -134 668
rect -128 653 -126 656
rect -76 653 -74 668
rect -68 653 -66 656
rect 221 689 232 691
rect 272 689 287 691
rect 327 689 331 691
rect 221 681 232 683
rect 272 681 287 683
rect 327 681 331 683
rect -325 613 -323 616
rect -445 605 -443 609
rect -437 605 -435 609
rect -385 605 -383 609
rect -377 605 -375 609
rect -16 640 -14 654
rect 387 652 398 654
rect 438 652 453 654
rect 493 652 497 654
rect 387 644 398 646
rect 438 644 453 646
rect 493 644 497 646
rect 65 624 76 626
rect 116 624 131 626
rect 171 624 175 626
rect -16 617 -14 620
rect 65 616 76 618
rect 116 616 131 618
rect 171 616 175 618
rect -136 609 -134 613
rect -128 609 -126 613
rect -76 609 -74 613
rect -68 609 -66 613
rect 221 603 232 605
rect 272 603 287 605
rect 327 603 331 605
rect -188 595 -186 599
rect -497 591 -495 595
rect 221 595 232 597
rect 272 595 287 597
rect 327 595 331 597
rect 596 579 598 582
rect 596 525 598 539
rect 193 514 204 516
rect 244 514 259 516
rect 299 514 303 516
rect 193 506 204 508
rect 244 506 259 508
rect 299 506 303 508
rect 596 502 598 505
rect 908 423 919 425
rect 959 423 983 425
rect 1063 423 1066 425
rect 908 415 919 417
rect 959 415 983 417
rect 1063 415 1066 417
rect -578 400 -576 413
rect -570 400 -568 413
rect -240 400 -238 413
rect -232 400 -230 413
rect 215 407 226 409
rect 266 407 281 409
rect 321 407 325 409
rect -526 373 -524 384
rect -466 373 -464 384
rect -406 359 -404 362
rect -578 284 -576 320
rect -570 309 -568 320
rect -526 318 -524 333
rect -518 318 -516 321
rect -466 318 -464 333
rect -458 318 -456 321
rect 908 407 919 409
rect 959 407 983 409
rect 1063 407 1066 409
rect 215 399 226 401
rect 266 399 281 401
rect 321 399 325 401
rect 908 399 919 401
rect 959 399 983 401
rect 1063 399 1066 401
rect 908 391 919 393
rect 959 391 983 393
rect 1063 391 1066 393
rect -188 373 -186 384
rect -128 373 -126 384
rect 381 370 392 372
rect 432 370 447 372
rect 487 370 491 372
rect -68 359 -66 362
rect 381 362 392 364
rect 432 362 447 364
rect 487 362 491 364
rect -406 305 -404 319
rect -406 282 -404 285
rect -240 284 -238 320
rect -232 309 -230 320
rect -188 318 -186 333
rect -180 318 -178 321
rect -128 318 -126 333
rect -120 318 -118 321
rect 1629 348 1631 361
rect 1637 348 1639 361
rect 59 342 70 344
rect 110 342 125 344
rect 165 342 169 344
rect 1192 338 1203 340
rect 1243 338 1267 340
rect 1347 338 1350 340
rect 59 334 70 336
rect 110 334 125 336
rect 165 334 169 336
rect 1192 330 1203 332
rect 1243 330 1267 332
rect 1347 330 1350 332
rect 215 321 226 323
rect 266 321 281 323
rect 321 321 325 323
rect 1192 322 1203 324
rect 1243 322 1267 324
rect 1347 322 1350 324
rect -526 274 -524 278
rect -518 274 -516 278
rect -466 274 -464 278
rect -458 274 -456 278
rect -68 305 -66 319
rect 215 313 226 315
rect 266 313 281 315
rect 321 313 325 315
rect 1192 314 1203 316
rect 1243 314 1267 316
rect 1347 314 1350 316
rect 1192 306 1203 308
rect 1243 306 1267 308
rect 1347 306 1350 308
rect -68 282 -66 285
rect -188 274 -186 278
rect -180 274 -178 278
rect -128 274 -126 278
rect -120 274 -118 278
rect -578 260 -576 264
rect -240 260 -238 264
rect 1681 321 1683 332
rect 1741 321 1743 332
rect 1801 307 1803 310
rect 930 262 941 264
rect 981 262 1005 264
rect 1085 262 1088 264
rect 930 254 941 256
rect 981 254 1005 256
rect 1085 254 1088 256
rect 930 246 941 248
rect 981 246 1005 248
rect 1085 246 1088 248
rect 930 238 941 240
rect 981 238 1005 240
rect 1085 238 1088 240
rect 187 232 198 234
rect 238 232 253 234
rect 293 232 297 234
rect 1629 232 1631 268
rect 1637 257 1639 268
rect 1681 266 1683 281
rect 1689 266 1691 269
rect 1741 266 1743 281
rect 1749 266 1751 269
rect 187 224 198 226
rect 238 224 253 226
rect 293 224 297 226
rect 1801 253 1803 267
rect 1801 230 1803 233
rect 1681 222 1683 226
rect 1689 222 1691 226
rect 1741 222 1743 226
rect 1749 222 1751 226
rect 1629 208 1631 212
rect 943 118 954 120
rect 994 118 1012 120
rect 1072 118 1077 120
rect 943 110 954 112
rect 994 110 1012 112
rect 1072 110 1077 112
rect 943 102 954 104
rect 994 102 1012 104
rect 1072 102 1077 104
rect 963 28 974 30
rect 1014 28 1029 30
rect 1069 28 1073 30
rect 963 20 974 22
rect 1014 20 1029 22
rect 1069 20 1073 22
<< polycontact >>
rect -120 1877 -116 1881
rect -112 1877 -108 1881
rect 682 1865 686 1869
rect 690 1865 694 1869
rect -68 1848 -64 1852
rect -8 1848 -4 1852
rect -60 1785 -56 1789
rect 0 1785 4 1789
rect 49 1772 53 1776
rect 734 1836 738 1840
rect 794 1836 798 1840
rect 742 1773 746 1777
rect 802 1773 806 1777
rect 241 1722 245 1726
rect 241 1714 245 1718
rect 851 1760 855 1764
rect 2180 1726 2184 1730
rect 2188 1726 2192 1730
rect 407 1685 411 1689
rect 407 1677 411 1681
rect 85 1657 89 1661
rect 85 1649 89 1653
rect 241 1636 245 1640
rect -190 1627 -186 1631
rect -182 1627 -178 1631
rect 241 1628 245 1632
rect 1749 1636 1753 1640
rect 1749 1628 1753 1632
rect 2232 1697 2236 1701
rect 2292 1697 2296 1701
rect -138 1598 -134 1602
rect -78 1598 -74 1602
rect 1915 1599 1919 1603
rect 1915 1591 1919 1595
rect 2240 1634 2244 1638
rect 2300 1634 2304 1638
rect -130 1535 -126 1539
rect -70 1535 -66 1539
rect 616 1562 620 1566
rect 1593 1571 1597 1575
rect 2349 1621 2353 1625
rect 1593 1563 1597 1567
rect 213 1547 217 1551
rect 213 1539 217 1543
rect 1749 1550 1753 1554
rect 1749 1542 1753 1546
rect -21 1522 -17 1526
rect 2184 1466 2188 1470
rect 2192 1466 2196 1470
rect -515 1400 -511 1404
rect -507 1400 -503 1404
rect -158 1403 -154 1407
rect -150 1403 -146 1407
rect -463 1371 -459 1375
rect -403 1371 -399 1375
rect -455 1308 -451 1312
rect -395 1308 -391 1312
rect -106 1374 -102 1378
rect -46 1374 -42 1378
rect 248 1371 252 1375
rect 2236 1437 2240 1441
rect 2296 1437 2300 1441
rect 248 1363 252 1367
rect 1749 1361 1753 1365
rect 1749 1353 1753 1357
rect -346 1295 -342 1299
rect -98 1311 -94 1315
rect -38 1311 -34 1315
rect 414 1334 418 1338
rect 2244 1374 2248 1378
rect 2304 1374 2308 1378
rect 414 1326 418 1330
rect 1915 1324 1919 1328
rect 1915 1316 1919 1320
rect 2353 1361 2357 1365
rect 11 1298 15 1302
rect 92 1306 96 1310
rect 92 1298 96 1302
rect 956 1301 960 1305
rect 956 1293 960 1297
rect 1593 1296 1597 1300
rect 248 1285 252 1289
rect 1593 1288 1597 1292
rect 248 1277 252 1281
rect 1749 1275 1753 1279
rect 1749 1267 1753 1271
rect 1180 1236 1184 1240
rect 2192 1242 2196 1246
rect 2200 1242 2204 1246
rect 1180 1228 1184 1232
rect 619 1211 623 1215
rect 220 1196 224 1200
rect 220 1188 224 1192
rect 1751 1167 1755 1171
rect 1751 1159 1755 1163
rect 2244 1213 2248 1217
rect 2304 1213 2308 1217
rect 1917 1130 1921 1134
rect 1917 1122 1921 1126
rect 2252 1150 2256 1154
rect 2312 1150 2316 1154
rect 1595 1102 1599 1106
rect -208 1096 -204 1100
rect -200 1096 -196 1100
rect -539 1086 -535 1090
rect -531 1086 -527 1090
rect 950 1094 954 1098
rect 950 1086 954 1090
rect 1595 1094 1599 1098
rect 2361 1137 2365 1141
rect -487 1057 -483 1061
rect -427 1057 -423 1061
rect -479 994 -475 998
rect -419 994 -415 998
rect 950 1078 954 1082
rect 1751 1081 1755 1085
rect 1751 1073 1755 1077
rect -156 1067 -152 1071
rect -96 1067 -92 1071
rect 1139 1053 1143 1057
rect 1139 1045 1143 1049
rect -370 981 -366 985
rect -148 1004 -144 1008
rect -88 1004 -84 1008
rect 218 1030 222 1034
rect 1139 1037 1143 1041
rect 218 1022 222 1026
rect 2185 1022 2189 1026
rect 2193 1022 2197 1026
rect 959 1010 963 1014
rect 959 1002 963 1006
rect -39 991 -35 995
rect 384 993 388 997
rect 384 985 388 989
rect 62 965 66 969
rect 1758 966 1762 970
rect 62 957 66 961
rect 1758 958 1762 962
rect 218 944 222 948
rect 218 936 222 940
rect 936 928 940 932
rect 1924 929 1928 933
rect 936 920 940 924
rect 1924 921 1928 925
rect 2237 993 2241 997
rect 2297 993 2301 997
rect 936 912 940 916
rect 936 904 940 908
rect 1602 901 1606 905
rect 1602 893 1606 897
rect 2245 930 2249 934
rect 2305 930 2309 934
rect 598 870 602 874
rect 1155 879 1159 883
rect 1758 880 1762 884
rect 1155 871 1159 875
rect 1758 872 1762 876
rect 2354 917 2358 921
rect 190 855 194 859
rect 190 847 194 851
rect 1155 863 1159 867
rect 1155 855 1159 859
rect 946 831 950 835
rect 946 823 950 827
rect 946 815 950 819
rect 955 758 959 762
rect -189 748 -185 752
rect -181 748 -177 752
rect 955 750 959 754
rect -498 744 -494 748
rect -490 744 -486 748
rect -446 715 -442 719
rect -386 715 -382 719
rect -438 652 -434 656
rect -378 652 -374 656
rect -137 719 -133 723
rect -77 719 -73 723
rect -329 639 -325 643
rect -129 656 -125 660
rect -69 656 -65 660
rect 217 688 221 692
rect 217 680 221 684
rect -20 643 -16 647
rect 383 651 387 655
rect 383 643 387 647
rect 61 623 65 627
rect 61 615 65 619
rect 217 602 221 606
rect 217 594 221 598
rect 592 528 596 532
rect 189 513 193 517
rect 189 505 193 509
rect 904 422 908 426
rect -579 413 -575 417
rect -571 413 -567 417
rect -241 413 -237 417
rect -233 413 -229 417
rect 904 414 908 418
rect 211 406 215 410
rect -527 384 -523 388
rect -467 384 -463 388
rect -519 321 -515 325
rect -459 321 -455 325
rect 211 398 215 402
rect 904 406 908 410
rect 904 398 908 402
rect 904 390 908 394
rect -189 384 -185 388
rect -129 384 -125 388
rect 377 369 381 373
rect 377 361 381 365
rect -410 308 -406 312
rect -181 321 -177 325
rect -121 321 -117 325
rect 1628 361 1632 365
rect 1636 361 1640 365
rect 55 341 59 345
rect 55 333 59 337
rect 1188 337 1192 341
rect 1188 329 1192 333
rect 211 320 215 324
rect 1188 321 1192 325
rect -72 308 -68 312
rect 211 312 215 316
rect 1188 313 1192 317
rect 1188 305 1192 309
rect 926 261 930 265
rect 1680 332 1684 336
rect 1740 332 1744 336
rect 926 253 930 257
rect 926 245 930 249
rect 183 231 187 235
rect 926 237 930 241
rect 1688 269 1692 273
rect 1748 269 1752 273
rect 183 223 187 227
rect 1797 256 1801 260
rect 939 117 943 121
rect 939 109 943 113
rect 939 101 943 105
rect 959 27 963 31
rect 959 19 963 23
<< metal1 >>
rect -78 1902 47 1906
rect -78 1894 -74 1902
rect -135 1890 -78 1894
rect -152 1883 -144 1887
rect -135 1869 -131 1890
rect -122 1882 -116 1887
rect -120 1881 -116 1882
rect -112 1881 -64 1884
rect -93 1870 -89 1881
rect -135 1865 -120 1869
rect -124 1864 -120 1865
rect -68 1857 -64 1881
rect -68 1852 -27 1857
rect -78 1843 -73 1847
rect -78 1838 -68 1843
rect -72 1837 -68 1838
rect -39 1801 -35 1806
rect -60 1797 -35 1801
rect -108 1768 -104 1784
rect -89 1785 -60 1789
rect -89 1768 -85 1785
rect -116 1764 -85 1768
rect -116 1748 -112 1764
rect -39 1742 -35 1797
rect -32 1790 -27 1852
rect -21 1841 -17 1902
rect 41 1900 47 1902
rect 41 1896 54 1900
rect -9 1852 -4 1856
rect -21 1837 -8 1841
rect 41 1831 47 1896
rect 724 1890 849 1894
rect 724 1882 728 1890
rect 667 1878 724 1882
rect 643 1873 658 1875
rect 573 1871 658 1873
rect 573 1869 647 1871
rect 41 1827 52 1831
rect 48 1823 52 1827
rect -4 1793 35 1797
rect -32 1789 4 1790
rect -32 1785 0 1789
rect -72 1732 -68 1742
rect -56 1738 -35 1742
rect 31 1775 35 1793
rect 41 1775 49 1776
rect -124 1725 -120 1728
rect -72 1727 -66 1732
rect -126 1720 -120 1725
rect -126 1710 -121 1720
rect -132 1707 -121 1710
rect -71 1708 -66 1727
rect -12 1708 -8 1742
rect 4 1730 8 1742
rect 25 1772 49 1775
rect 56 1775 60 1783
rect 25 1770 43 1772
rect 56 1771 72 1775
rect 25 1730 30 1770
rect 56 1769 60 1771
rect 48 1740 52 1749
rect 4 1725 30 1730
rect 43 1736 52 1740
rect 43 1708 48 1736
rect -71 1707 48 1708
rect -132 1706 48 1707
rect -126 1703 48 1706
rect -126 1702 -66 1703
rect 68 1661 72 1771
rect 304 1740 308 1741
rect 304 1736 406 1740
rect 304 1730 308 1736
rect 249 1726 256 1730
rect 304 1726 311 1730
rect 237 1725 241 1726
rect 81 1722 241 1725
rect 81 1721 240 1722
rect 81 1661 85 1721
rect 148 1714 241 1718
rect 249 1714 253 1726
rect 304 1722 308 1726
rect 296 1718 308 1722
rect 148 1678 152 1714
rect 249 1710 256 1714
rect 351 1710 362 1714
rect 244 1706 253 1710
rect 244 1702 248 1706
rect 402 1689 406 1736
rect 573 1707 577 1869
rect 667 1857 671 1878
rect 680 1870 686 1875
rect 682 1869 686 1870
rect 690 1869 738 1872
rect 709 1861 713 1869
rect 667 1853 682 1857
rect 678 1852 682 1853
rect 734 1845 738 1869
rect 734 1840 775 1845
rect 724 1831 729 1835
rect 724 1826 734 1831
rect 730 1825 734 1826
rect 763 1789 767 1794
rect 742 1785 767 1789
rect 694 1756 698 1772
rect 713 1773 742 1777
rect 713 1756 717 1773
rect 686 1752 717 1756
rect 686 1736 690 1752
rect 763 1730 767 1785
rect 770 1778 775 1840
rect 781 1829 785 1890
rect 843 1888 849 1890
rect 843 1884 856 1888
rect 793 1840 798 1844
rect 781 1825 794 1829
rect 843 1819 849 1884
rect 843 1815 854 1819
rect 850 1811 854 1815
rect 798 1781 837 1785
rect 770 1777 806 1778
rect 770 1773 802 1777
rect 730 1720 734 1730
rect 746 1726 767 1730
rect 833 1763 837 1781
rect 843 1763 851 1764
rect 678 1713 682 1716
rect 730 1715 736 1720
rect 470 1703 577 1707
rect 676 1708 682 1713
rect 470 1693 474 1703
rect 676 1698 681 1708
rect 670 1695 681 1698
rect 731 1696 736 1715
rect 790 1696 794 1730
rect 806 1718 810 1730
rect 827 1760 851 1763
rect 858 1763 862 1771
rect 827 1758 845 1760
rect 858 1759 868 1763
rect 827 1718 832 1758
rect 858 1757 862 1759
rect 2222 1752 2347 1755
rect 2222 1751 2354 1752
rect 2222 1743 2226 1751
rect 2165 1739 2222 1743
rect 850 1728 854 1737
rect 806 1713 832 1718
rect 845 1724 854 1728
rect 1978 1731 2156 1735
rect 845 1696 850 1724
rect 731 1695 850 1696
rect 670 1694 850 1695
rect 415 1689 422 1693
rect 470 1689 477 1693
rect 676 1691 850 1694
rect 676 1690 736 1691
rect 402 1685 407 1689
rect 403 1679 407 1681
rect 148 1674 239 1678
rect 148 1665 152 1674
rect 93 1661 100 1665
rect 148 1661 155 1665
rect 31 1657 52 1661
rect 57 1657 85 1661
rect -148 1652 -23 1656
rect -148 1644 -144 1652
rect -205 1640 -148 1644
rect -221 1633 -214 1637
rect -205 1619 -201 1640
rect -192 1632 -186 1637
rect -190 1631 -186 1632
rect -182 1631 -134 1634
rect -163 1620 -159 1631
rect -205 1615 -190 1619
rect -194 1614 -190 1615
rect -138 1607 -134 1631
rect -138 1602 -97 1607
rect -148 1593 -143 1597
rect -148 1588 -138 1593
rect -142 1587 -138 1588
rect -109 1551 -105 1556
rect -130 1547 -105 1551
rect -178 1518 -174 1534
rect -159 1535 -130 1539
rect -159 1518 -155 1535
rect -186 1514 -155 1518
rect -186 1498 -182 1514
rect -109 1492 -105 1547
rect -102 1540 -97 1602
rect -91 1591 -87 1652
rect -29 1650 -23 1652
rect -29 1646 -16 1650
rect -79 1602 -74 1606
rect -91 1587 -78 1591
rect -29 1581 -23 1646
rect 37 1649 85 1653
rect 93 1649 97 1661
rect 148 1657 152 1661
rect 140 1653 152 1657
rect 37 1643 41 1649
rect 31 1639 41 1643
rect -29 1577 -18 1581
rect -22 1573 -18 1577
rect -74 1543 -35 1547
rect -102 1539 -66 1540
rect -102 1535 -70 1539
rect -142 1482 -138 1492
rect -126 1488 -105 1492
rect -39 1525 -35 1543
rect -29 1525 -21 1526
rect -194 1475 -190 1478
rect -142 1477 -136 1482
rect -196 1470 -190 1475
rect -196 1460 -191 1470
rect -202 1457 -191 1460
rect -141 1458 -136 1477
rect -82 1458 -78 1492
rect -66 1480 -62 1492
rect -45 1522 -21 1525
rect -14 1525 -10 1533
rect 33 1525 37 1639
rect 65 1615 69 1649
rect 93 1645 100 1649
rect 195 1645 206 1649
rect 88 1641 97 1645
rect 88 1637 92 1641
rect 235 1640 239 1674
rect 304 1675 407 1679
rect 415 1677 419 1689
rect 470 1685 474 1689
rect 462 1681 474 1685
rect 304 1644 308 1675
rect 415 1673 422 1677
rect 517 1673 528 1677
rect 410 1669 419 1673
rect 410 1665 414 1669
rect 1812 1654 1816 1655
rect 1812 1650 1914 1654
rect 1812 1644 1816 1650
rect 249 1640 256 1644
rect 304 1640 311 1644
rect 1757 1640 1764 1644
rect 1812 1640 1819 1644
rect 235 1636 241 1640
rect 237 1630 241 1632
rect 155 1628 241 1630
rect 249 1628 253 1640
rect 304 1636 308 1640
rect 1745 1639 1749 1640
rect 1589 1636 1749 1639
rect 296 1632 308 1636
rect 1589 1635 1748 1636
rect 155 1626 240 1628
rect 155 1615 159 1626
rect 65 1611 159 1615
rect 200 1551 204 1626
rect 249 1624 256 1628
rect 351 1624 362 1628
rect 244 1620 253 1624
rect 244 1616 248 1620
rect 611 1619 633 1623
rect 615 1613 619 1619
rect 1589 1580 1593 1635
rect 1527 1576 1593 1580
rect 1656 1628 1749 1632
rect 1757 1628 1761 1640
rect 1812 1636 1816 1640
rect 1804 1632 1816 1636
rect 1656 1592 1660 1628
rect 1757 1624 1764 1628
rect 1859 1624 1870 1628
rect 1752 1620 1761 1624
rect 1752 1616 1756 1620
rect 1910 1603 1914 1650
rect 1978 1607 1982 1731
rect 2165 1718 2169 1739
rect 2178 1731 2184 1736
rect 2180 1730 2184 1731
rect 2188 1730 2204 1733
rect 2210 1730 2236 1733
rect 2165 1714 2180 1718
rect 2176 1713 2180 1714
rect 2232 1706 2236 1730
rect 2232 1701 2273 1706
rect 2222 1692 2227 1696
rect 2222 1687 2232 1692
rect 2228 1686 2232 1687
rect 2261 1650 2265 1655
rect 2240 1646 2265 1650
rect 2192 1617 2196 1633
rect 2211 1634 2240 1638
rect 2211 1617 2215 1634
rect 2184 1613 2215 1617
rect 1923 1603 1930 1607
rect 1978 1603 1985 1607
rect 1910 1599 1915 1603
rect 1911 1593 1915 1595
rect 1656 1588 1747 1592
rect 1656 1579 1660 1588
rect 623 1566 627 1573
rect 1589 1571 1593 1576
rect 1601 1575 1608 1579
rect 1656 1575 1663 1579
rect 1568 1567 1579 1568
rect 276 1562 616 1566
rect 623 1565 641 1566
rect 1568 1565 1593 1567
rect 623 1563 1593 1565
rect 1601 1563 1605 1575
rect 1656 1571 1660 1575
rect 1648 1567 1660 1571
rect 623 1562 1579 1563
rect 276 1555 280 1562
rect 623 1559 627 1562
rect 221 1551 228 1555
rect 276 1551 283 1555
rect 200 1547 213 1551
rect 212 1539 213 1543
rect 221 1539 225 1551
rect 276 1547 280 1551
rect 268 1543 280 1547
rect 221 1535 228 1539
rect 323 1535 332 1539
rect 637 1561 1579 1562
rect 216 1531 225 1535
rect 615 1535 619 1539
rect 609 1531 633 1535
rect 216 1528 220 1531
rect -45 1520 -27 1522
rect -14 1521 37 1525
rect -45 1480 -40 1520
rect -14 1519 -10 1521
rect -22 1490 -18 1499
rect -66 1475 -40 1480
rect -27 1486 -18 1490
rect -27 1458 -22 1486
rect -141 1457 -22 1458
rect -202 1456 -22 1457
rect -196 1453 -22 1456
rect -196 1452 -136 1453
rect -473 1425 -348 1429
rect -473 1417 -469 1425
rect -530 1413 -473 1417
rect -554 1408 -539 1410
rect -564 1406 -539 1408
rect -564 1404 -550 1406
rect -530 1392 -526 1413
rect -517 1405 -511 1410
rect -515 1404 -511 1405
rect -507 1404 -459 1407
rect -488 1393 -484 1404
rect -530 1388 -515 1392
rect -519 1387 -515 1388
rect -463 1380 -459 1404
rect -463 1375 -422 1380
rect -473 1366 -468 1370
rect -473 1361 -463 1366
rect -467 1360 -463 1361
rect -434 1324 -430 1329
rect -455 1320 -430 1324
rect -503 1291 -499 1307
rect -484 1308 -455 1312
rect -484 1291 -480 1308
rect -511 1287 -480 1291
rect -511 1271 -507 1287
rect -434 1265 -430 1320
rect -427 1313 -422 1375
rect -416 1364 -412 1425
rect -354 1423 -348 1425
rect -116 1428 9 1432
rect -354 1419 -341 1423
rect -404 1375 -399 1379
rect -416 1360 -403 1364
rect -354 1354 -348 1419
rect -116 1420 -112 1428
rect -173 1416 -116 1420
rect -197 1411 -182 1413
rect -207 1409 -182 1411
rect -207 1407 -193 1409
rect -173 1395 -169 1416
rect -160 1408 -154 1413
rect -158 1407 -154 1408
rect -150 1407 -102 1410
rect -131 1396 -127 1407
rect -173 1391 -158 1395
rect -162 1390 -158 1391
rect -354 1350 -343 1354
rect -347 1346 -343 1350
rect -399 1316 -360 1320
rect -427 1312 -391 1313
rect -427 1308 -395 1312
rect -467 1255 -463 1265
rect -451 1261 -430 1265
rect -364 1298 -360 1316
rect -106 1383 -102 1407
rect -106 1378 -65 1383
rect -116 1369 -111 1373
rect -116 1364 -106 1369
rect -110 1363 -106 1364
rect -77 1327 -73 1332
rect -98 1323 -73 1327
rect -354 1298 -346 1299
rect -519 1248 -515 1251
rect -467 1250 -461 1255
rect -521 1243 -515 1248
rect -521 1233 -516 1243
rect -527 1230 -516 1233
rect -466 1231 -461 1250
rect -407 1231 -403 1265
rect -391 1253 -387 1265
rect -370 1295 -346 1298
rect -339 1298 -335 1306
rect -370 1293 -352 1295
rect -339 1294 -304 1298
rect -146 1294 -142 1310
rect -127 1311 -98 1315
rect -127 1294 -123 1311
rect -370 1253 -365 1293
rect -339 1292 -335 1294
rect -347 1263 -343 1272
rect -391 1248 -365 1253
rect -352 1259 -343 1263
rect -352 1231 -347 1259
rect -466 1230 -347 1231
rect -527 1229 -347 1230
rect -521 1226 -347 1229
rect -521 1225 -461 1226
rect -308 1205 -304 1294
rect -154 1290 -123 1294
rect -154 1274 -150 1290
rect -77 1268 -73 1323
rect -70 1316 -65 1378
rect -59 1367 -55 1428
rect 3 1426 9 1428
rect 3 1422 16 1426
rect -47 1378 -42 1382
rect -59 1363 -46 1367
rect 3 1357 9 1422
rect 311 1389 315 1390
rect 311 1385 413 1389
rect 311 1379 315 1385
rect 256 1375 263 1379
rect 311 1375 318 1379
rect 244 1374 248 1375
rect 88 1371 248 1374
rect 88 1370 247 1371
rect 3 1353 14 1357
rect 10 1349 14 1353
rect -42 1319 -3 1323
rect -70 1315 -34 1316
rect -70 1311 -38 1315
rect -110 1258 -106 1268
rect -94 1264 -73 1268
rect -7 1301 -3 1319
rect 88 1310 92 1370
rect 155 1363 248 1367
rect 256 1363 260 1375
rect 311 1371 315 1375
rect 303 1367 315 1371
rect 155 1327 159 1363
rect 256 1359 263 1363
rect 358 1359 369 1363
rect 251 1355 260 1359
rect 251 1351 255 1355
rect 409 1338 413 1385
rect 477 1352 601 1356
rect 477 1342 481 1352
rect 422 1338 429 1342
rect 477 1338 484 1342
rect 409 1334 414 1338
rect 410 1328 414 1330
rect 155 1323 246 1327
rect 155 1314 159 1323
rect 100 1310 107 1314
rect 155 1310 162 1314
rect 3 1301 11 1302
rect -162 1251 -158 1254
rect -110 1253 -104 1258
rect -164 1246 -158 1251
rect -164 1236 -159 1246
rect -170 1233 -159 1236
rect -109 1234 -104 1253
rect -50 1234 -46 1268
rect -34 1256 -30 1268
rect -13 1298 11 1301
rect 18 1301 22 1309
rect 31 1306 59 1310
rect 31 1301 35 1306
rect 64 1306 92 1310
rect -13 1296 5 1298
rect 18 1297 35 1301
rect 44 1298 92 1302
rect 100 1298 104 1310
rect 155 1306 159 1310
rect 147 1302 159 1306
rect -13 1256 -8 1296
rect 18 1295 22 1297
rect 44 1292 48 1298
rect 38 1288 48 1292
rect 10 1266 14 1275
rect -34 1251 -8 1256
rect 5 1262 14 1266
rect 5 1234 10 1262
rect -109 1233 10 1234
rect -170 1232 10 1233
rect -164 1229 10 1232
rect -164 1228 -104 1229
rect 38 1225 42 1288
rect 72 1264 76 1298
rect 100 1294 107 1298
rect 202 1294 213 1298
rect 95 1290 104 1294
rect 95 1286 99 1290
rect 242 1289 246 1323
rect 311 1324 414 1328
rect 422 1326 426 1338
rect 477 1334 481 1338
rect 469 1330 481 1334
rect 311 1293 315 1324
rect 422 1322 429 1326
rect 524 1322 535 1326
rect 417 1318 426 1322
rect 417 1314 421 1318
rect 587 1297 591 1352
rect 637 1307 641 1561
rect 1568 1557 1579 1561
rect 1601 1559 1608 1563
rect 1703 1559 1714 1563
rect 1573 1529 1577 1557
rect 1596 1555 1605 1559
rect 1596 1551 1600 1555
rect 1743 1554 1747 1588
rect 1812 1589 1915 1593
rect 1923 1591 1927 1603
rect 1978 1599 1982 1603
rect 1970 1595 1982 1599
rect 2184 1597 2188 1613
rect 1812 1558 1816 1589
rect 1923 1587 1930 1591
rect 2025 1587 2036 1591
rect 1918 1583 1927 1587
rect 1918 1579 1922 1583
rect 2261 1591 2265 1646
rect 2268 1639 2273 1701
rect 2279 1690 2283 1751
rect 2341 1748 2354 1751
rect 2291 1701 2296 1705
rect 2279 1686 2292 1690
rect 2341 1680 2347 1748
rect 2341 1676 2352 1680
rect 2348 1672 2352 1676
rect 2296 1642 2335 1646
rect 2268 1638 2304 1639
rect 2268 1634 2300 1638
rect 2228 1581 2232 1591
rect 2244 1587 2265 1591
rect 2331 1624 2335 1642
rect 2341 1624 2349 1625
rect 2176 1574 2180 1577
rect 2228 1576 2234 1581
rect 2174 1569 2180 1574
rect 1757 1554 1764 1558
rect 1812 1554 1819 1558
rect 2174 1557 2179 1569
rect 1743 1550 1749 1554
rect 1745 1544 1749 1546
rect 1663 1542 1749 1544
rect 1757 1542 1761 1554
rect 1812 1550 1816 1554
rect 2168 1556 2179 1557
rect 2229 1557 2234 1576
rect 2288 1557 2292 1591
rect 2304 1579 2308 1591
rect 2325 1621 2349 1624
rect 2356 1624 2360 1632
rect 2325 1619 2343 1621
rect 2356 1620 2366 1624
rect 2325 1579 2330 1619
rect 2356 1618 2360 1620
rect 2348 1589 2352 1598
rect 2304 1574 2330 1579
rect 2343 1585 2352 1589
rect 2343 1557 2348 1585
rect 2229 1556 2348 1557
rect 2168 1553 2348 1556
rect 2174 1552 2348 1553
rect 2174 1551 2234 1552
rect 1804 1546 1816 1550
rect 1663 1540 1748 1542
rect 1663 1529 1667 1540
rect 1757 1538 1764 1542
rect 1859 1538 1870 1542
rect 1752 1534 1761 1538
rect 1752 1530 1756 1534
rect 1573 1525 1667 1529
rect 2226 1492 2351 1495
rect 2226 1491 2358 1492
rect 2226 1483 2230 1491
rect 2169 1479 2226 1483
rect 1978 1471 2160 1475
rect 1812 1379 1816 1380
rect 1812 1375 1914 1379
rect 1812 1369 1816 1375
rect 1757 1365 1764 1369
rect 1812 1365 1819 1369
rect 1745 1364 1749 1365
rect 1589 1361 1749 1364
rect 1589 1360 1748 1361
rect 775 1307 779 1310
rect 1019 1312 1143 1316
rect 1019 1309 1023 1312
rect 637 1305 955 1307
rect 964 1305 971 1309
rect 1019 1305 1026 1309
rect 637 1303 923 1305
rect 928 1303 956 1305
rect 946 1301 956 1303
rect 946 1300 955 1301
rect 587 1293 956 1297
rect 964 1293 968 1305
rect 1019 1301 1023 1305
rect 1011 1297 1023 1301
rect 256 1289 263 1293
rect 311 1289 318 1293
rect 850 1290 854 1293
rect 932 1290 936 1293
rect 242 1285 248 1289
rect 244 1279 248 1281
rect 162 1277 248 1279
rect 256 1277 260 1289
rect 311 1285 315 1289
rect 964 1289 971 1293
rect 1066 1289 1075 1293
rect 959 1285 968 1289
rect 303 1281 315 1285
rect 959 1282 963 1285
rect 162 1275 247 1277
rect 162 1264 166 1275
rect 72 1260 166 1264
rect -158 1221 42 1225
rect -158 1205 -154 1221
rect -308 1201 -154 1205
rect 207 1200 211 1275
rect 256 1273 263 1277
rect 358 1273 369 1277
rect 251 1269 260 1273
rect 251 1265 255 1269
rect 614 1268 636 1272
rect 618 1262 622 1268
rect 1139 1240 1143 1312
rect 1589 1300 1593 1360
rect 1656 1353 1749 1357
rect 1757 1353 1761 1365
rect 1812 1361 1816 1365
rect 1804 1357 1816 1361
rect 1656 1317 1660 1353
rect 1757 1349 1764 1353
rect 1859 1349 1870 1353
rect 1752 1345 1761 1349
rect 1752 1341 1756 1345
rect 1910 1328 1914 1375
rect 1978 1332 1982 1471
rect 2169 1458 2173 1479
rect 2182 1471 2188 1476
rect 2184 1470 2188 1471
rect 2192 1470 2204 1473
rect 2210 1470 2240 1473
rect 2169 1454 2184 1458
rect 2180 1453 2184 1454
rect 2236 1446 2240 1470
rect 2236 1441 2277 1446
rect 2226 1432 2231 1436
rect 2226 1427 2236 1432
rect 2232 1426 2236 1427
rect 2265 1390 2269 1395
rect 2244 1386 2269 1390
rect 2196 1357 2200 1373
rect 2215 1374 2244 1378
rect 2215 1357 2219 1374
rect 2188 1353 2219 1357
rect 2188 1337 2192 1353
rect 1923 1328 1930 1332
rect 1978 1328 1985 1332
rect 1910 1324 1915 1328
rect 1911 1318 1915 1320
rect 1656 1313 1747 1317
rect 1656 1304 1660 1313
rect 1601 1300 1608 1304
rect 1656 1300 1663 1304
rect 1540 1296 1593 1300
rect 1540 1295 1592 1296
rect 1573 1291 1593 1292
rect 1487 1288 1593 1291
rect 1601 1288 1605 1300
rect 1656 1296 1660 1300
rect 1648 1292 1660 1296
rect 1487 1287 1578 1288
rect 1487 1268 1491 1287
rect 1243 1264 1491 1268
rect 1243 1244 1247 1264
rect 1188 1240 1195 1244
rect 1243 1240 1250 1244
rect 1139 1236 1180 1240
rect 626 1215 630 1222
rect 1139 1228 1180 1232
rect 1188 1228 1192 1240
rect 1243 1236 1247 1240
rect 1235 1232 1247 1236
rect 283 1211 619 1215
rect 626 1213 914 1215
rect 626 1211 862 1213
rect 283 1204 287 1211
rect 228 1200 235 1204
rect 283 1200 290 1204
rect 207 1196 220 1200
rect 219 1188 220 1192
rect 228 1188 232 1200
rect 283 1196 287 1200
rect 275 1192 287 1196
rect 228 1184 235 1188
rect 330 1184 339 1188
rect 223 1180 232 1184
rect 223 1177 227 1180
rect 564 1168 568 1211
rect 626 1208 630 1211
rect 684 1204 688 1211
rect 867 1211 914 1213
rect 618 1184 622 1188
rect 612 1180 636 1184
rect 656 1172 1001 1176
rect 1139 1168 1143 1228
rect 1188 1224 1195 1228
rect 1290 1224 1299 1228
rect 1183 1220 1192 1224
rect 1183 1217 1187 1220
rect 564 1164 1143 1168
rect -166 1121 -41 1125
rect -497 1111 -372 1115
rect -166 1113 -162 1121
rect -497 1103 -493 1111
rect -554 1099 -497 1103
rect -578 1094 -563 1096
rect -588 1092 -563 1094
rect -588 1090 -574 1092
rect -554 1078 -550 1099
rect -541 1091 -535 1096
rect -539 1090 -535 1091
rect -531 1090 -483 1093
rect -512 1079 -508 1090
rect -554 1074 -539 1078
rect -543 1073 -539 1074
rect -487 1066 -483 1090
rect -487 1061 -446 1066
rect -497 1052 -492 1056
rect -497 1047 -487 1052
rect -491 1046 -487 1047
rect -458 1010 -454 1015
rect -479 1006 -454 1010
rect -527 977 -523 993
rect -508 994 -479 998
rect -508 977 -504 994
rect -535 973 -504 977
rect -535 957 -531 973
rect -458 951 -454 1006
rect -451 999 -446 1061
rect -440 1050 -436 1111
rect -378 1109 -372 1111
rect -223 1109 -166 1113
rect -378 1105 -365 1109
rect -428 1061 -423 1065
rect -440 1046 -427 1050
rect -378 1040 -372 1105
rect -247 1104 -232 1106
rect -257 1102 -232 1104
rect -257 1100 -243 1102
rect -223 1088 -219 1109
rect -210 1101 -204 1106
rect -208 1100 -204 1101
rect -200 1100 -152 1103
rect -181 1089 -177 1100
rect -223 1084 -208 1088
rect -212 1083 -208 1084
rect -378 1036 -367 1040
rect -371 1032 -367 1036
rect -423 1002 -384 1006
rect -451 998 -415 999
rect -451 994 -419 998
rect -491 941 -487 951
rect -475 947 -454 951
rect -388 984 -384 1002
rect -156 1076 -152 1100
rect -156 1071 -115 1076
rect -166 1062 -161 1066
rect -166 1057 -156 1062
rect -160 1056 -156 1057
rect -127 1020 -123 1025
rect -148 1016 -123 1020
rect -378 984 -370 985
rect -543 934 -539 937
rect -491 936 -485 941
rect -545 929 -539 934
rect -545 919 -540 929
rect -551 916 -540 919
rect -490 917 -485 936
rect -431 917 -427 951
rect -415 939 -411 951
rect -394 981 -370 984
rect -363 984 -359 992
rect -196 987 -192 1003
rect -177 1004 -148 1008
rect -177 987 -173 1004
rect -394 979 -376 981
rect -363 980 -340 984
rect -394 939 -389 979
rect -363 978 -359 980
rect -371 949 -367 958
rect -415 934 -389 939
rect -376 945 -367 949
rect -376 917 -371 945
rect -490 916 -371 917
rect -551 915 -371 916
rect -545 912 -371 915
rect -545 911 -485 912
rect -344 899 -340 980
rect -204 983 -173 987
rect -204 967 -200 983
rect -127 961 -123 1016
rect -120 1009 -115 1071
rect -109 1060 -105 1121
rect -47 1119 -41 1121
rect -47 1115 -34 1119
rect -97 1071 -92 1075
rect -109 1056 -96 1060
rect -47 1050 -41 1115
rect -47 1046 -36 1050
rect -40 1042 -36 1046
rect 281 1048 285 1049
rect 281 1044 383 1048
rect -92 1012 -53 1016
rect -120 1008 -84 1009
rect -120 1004 -88 1008
rect -160 951 -156 961
rect -144 957 -123 961
rect -57 994 -53 1012
rect 281 1038 285 1044
rect 226 1034 233 1038
rect 281 1034 288 1038
rect 214 1033 218 1034
rect -47 994 -39 995
rect -212 944 -208 947
rect -160 946 -154 951
rect -214 939 -208 944
rect -214 929 -209 939
rect -220 926 -209 929
rect -159 927 -154 946
rect -100 927 -96 961
rect -84 949 -80 961
rect -63 991 -39 994
rect -32 994 -28 1002
rect 58 1030 218 1033
rect 58 1029 217 1030
rect -63 989 -45 991
rect -32 990 -18 994
rect -63 949 -58 989
rect -32 988 -28 990
rect -22 969 -18 990
rect 58 969 62 1029
rect 125 1022 218 1026
rect 226 1022 230 1034
rect 281 1030 285 1034
rect 273 1026 285 1030
rect 125 986 129 1022
rect 226 1018 233 1022
rect 328 1018 339 1022
rect 221 1014 230 1018
rect 221 1010 225 1014
rect 379 997 383 1044
rect 651 1015 655 1146
rect 923 1090 927 1149
rect 932 1098 936 1149
rect 1001 1146 1005 1150
rect 1535 1146 1539 1269
rect 1573 1254 1577 1287
rect 1601 1284 1608 1288
rect 1703 1284 1714 1288
rect 1596 1280 1605 1284
rect 1596 1276 1600 1280
rect 1743 1279 1747 1313
rect 1812 1314 1915 1318
rect 1923 1316 1927 1328
rect 1978 1324 1982 1328
rect 1970 1320 1982 1324
rect 2265 1331 2269 1386
rect 2272 1379 2277 1441
rect 2283 1430 2287 1491
rect 2345 1488 2358 1491
rect 2295 1441 2300 1445
rect 2283 1426 2296 1430
rect 2345 1420 2351 1488
rect 2345 1416 2356 1420
rect 2352 1412 2356 1416
rect 2300 1382 2339 1386
rect 2272 1378 2308 1379
rect 2272 1374 2304 1378
rect 2232 1321 2236 1331
rect 2248 1327 2269 1331
rect 2335 1364 2339 1382
rect 2345 1364 2353 1365
rect 1812 1283 1816 1314
rect 1923 1312 1930 1316
rect 2025 1312 2036 1316
rect 2180 1314 2184 1317
rect 2232 1316 2238 1321
rect 1918 1308 1927 1312
rect 2178 1309 2184 1314
rect 1918 1304 1922 1308
rect 2178 1300 2183 1309
rect 2174 1296 2183 1300
rect 2233 1297 2238 1316
rect 2292 1297 2296 1331
rect 2308 1319 2312 1331
rect 2329 1361 2353 1364
rect 2360 1364 2364 1372
rect 2329 1359 2347 1361
rect 2360 1360 2370 1364
rect 2329 1319 2334 1359
rect 2360 1358 2364 1360
rect 2352 1329 2356 1338
rect 2308 1314 2334 1319
rect 2347 1325 2356 1329
rect 2347 1297 2352 1325
rect 2233 1296 2352 1297
rect 2178 1292 2352 1296
rect 2178 1291 2238 1292
rect 1757 1279 1764 1283
rect 1812 1279 1819 1283
rect 1743 1275 1749 1279
rect 1745 1269 1749 1271
rect 1663 1267 1749 1269
rect 1757 1267 1761 1279
rect 1812 1275 1816 1279
rect 1804 1271 1816 1275
rect 1663 1265 1748 1267
rect 1663 1254 1667 1265
rect 1757 1263 1764 1267
rect 1859 1263 1870 1267
rect 2234 1267 2359 1271
rect 1752 1259 1761 1263
rect 2234 1259 2238 1267
rect 1752 1255 1756 1259
rect 1573 1250 1667 1254
rect 2177 1255 2234 1259
rect 1980 1252 2172 1253
rect 1980 1249 2168 1252
rect 1814 1185 1818 1186
rect 1814 1181 1916 1185
rect 1814 1175 1818 1181
rect 1759 1171 1766 1175
rect 1814 1171 1821 1175
rect 1747 1170 1751 1171
rect 1001 1142 1539 1146
rect 1591 1167 1751 1170
rect 1591 1166 1750 1167
rect 1207 1105 1493 1109
rect 1005 1098 1023 1102
rect 932 1094 950 1098
rect 958 1090 965 1094
rect 923 1086 950 1090
rect 899 1078 950 1082
rect 958 1078 962 1090
rect 1009 1086 1013 1098
rect 1005 1082 1013 1086
rect 899 1015 903 1078
rect 958 1074 965 1078
rect 958 1068 962 1074
rect 1009 1057 1013 1082
rect 1083 1074 1100 1078
rect 1207 1061 1211 1105
rect 1489 1098 1493 1105
rect 1591 1108 1595 1166
rect 1658 1159 1751 1163
rect 1759 1159 1763 1171
rect 1814 1167 1818 1171
rect 1806 1163 1818 1167
rect 1658 1123 1662 1159
rect 1759 1155 1766 1159
rect 1861 1155 1872 1159
rect 1754 1151 1763 1155
rect 1754 1147 1758 1151
rect 1912 1134 1916 1181
rect 1980 1138 1984 1249
rect 2177 1234 2181 1255
rect 2190 1247 2196 1252
rect 2192 1246 2196 1247
rect 2200 1246 2214 1249
rect 2220 1246 2248 1249
rect 2177 1230 2192 1234
rect 2188 1229 2192 1230
rect 2244 1222 2248 1246
rect 2244 1217 2285 1222
rect 2234 1208 2239 1212
rect 2234 1203 2244 1208
rect 2240 1202 2244 1203
rect 2273 1166 2277 1171
rect 2252 1162 2277 1166
rect 1925 1134 1932 1138
rect 1980 1134 1987 1138
rect 1912 1130 1917 1134
rect 1913 1124 1917 1126
rect 1658 1119 1749 1123
rect 1658 1110 1662 1119
rect 1559 1104 1595 1108
rect 1603 1106 1610 1110
rect 1658 1106 1665 1110
rect 1591 1102 1595 1104
rect 1489 1094 1595 1098
rect 1603 1094 1607 1106
rect 1658 1102 1662 1106
rect 1650 1098 1662 1102
rect 1194 1057 1212 1061
rect 1575 1060 1579 1094
rect 1603 1090 1610 1094
rect 1705 1090 1716 1094
rect 1598 1086 1607 1090
rect 1598 1082 1602 1086
rect 1745 1085 1749 1119
rect 1814 1120 1917 1124
rect 1925 1122 1929 1134
rect 1980 1130 1984 1134
rect 2204 1133 2208 1149
rect 2223 1150 2252 1154
rect 2223 1133 2227 1150
rect 1972 1126 1984 1130
rect 2196 1129 2227 1133
rect 1814 1089 1818 1120
rect 1925 1118 1932 1122
rect 2027 1118 2038 1122
rect 1920 1114 1929 1118
rect 1920 1110 1924 1114
rect 2196 1113 2200 1129
rect 2273 1107 2277 1162
rect 2280 1155 2285 1217
rect 2291 1206 2295 1267
rect 2353 1259 2359 1267
rect 2353 1255 2366 1259
rect 2303 1217 2308 1221
rect 2291 1202 2304 1206
rect 2353 1196 2359 1255
rect 2353 1192 2364 1196
rect 2360 1188 2364 1192
rect 2308 1158 2347 1162
rect 2280 1154 2316 1155
rect 2280 1150 2312 1154
rect 2240 1097 2244 1107
rect 2256 1103 2277 1107
rect 2343 1140 2347 1158
rect 2353 1140 2361 1141
rect 2188 1090 2192 1093
rect 2240 1092 2246 1097
rect 1759 1085 1766 1089
rect 1814 1085 1821 1089
rect 2186 1085 2192 1090
rect 1745 1081 1751 1085
rect 1747 1075 1751 1077
rect 1665 1073 1751 1075
rect 1759 1073 1763 1085
rect 1814 1081 1818 1085
rect 1806 1077 1818 1081
rect 2186 1077 2191 1085
rect 1665 1071 1750 1073
rect 1665 1060 1669 1071
rect 1759 1069 1766 1073
rect 1861 1069 1872 1073
rect 2180 1073 2191 1077
rect 2186 1072 2191 1073
rect 2241 1073 2246 1092
rect 2300 1073 2304 1107
rect 2316 1095 2320 1107
rect 2337 1137 2361 1140
rect 2368 1140 2372 1148
rect 2337 1135 2355 1137
rect 2368 1136 2378 1140
rect 2337 1095 2342 1135
rect 2368 1134 2372 1136
rect 2360 1105 2364 1114
rect 2316 1090 2342 1095
rect 2355 1101 2364 1105
rect 2355 1073 2360 1101
rect 2241 1072 2360 1073
rect 1754 1065 1763 1069
rect 2186 1068 2360 1072
rect 2186 1067 2246 1068
rect 1754 1061 1758 1065
rect 1009 1053 1139 1057
rect 1147 1049 1154 1053
rect 1022 1045 1139 1049
rect 1022 1018 1026 1045
rect 1103 1037 1139 1041
rect 1147 1037 1151 1049
rect 1198 1045 1202 1057
rect 1575 1056 1669 1060
rect 2227 1047 2352 1051
rect 1194 1041 1202 1045
rect 2227 1039 2231 1047
rect 1147 1033 1154 1037
rect 1272 1033 1289 1037
rect 2170 1035 2227 1039
rect 1147 1027 1151 1033
rect 1987 1032 2165 1034
rect 1987 1030 2161 1032
rect 447 1014 945 1015
rect 967 1014 974 1018
rect 1022 1014 1029 1018
rect 447 1011 959 1014
rect 447 1001 451 1011
rect 725 1010 734 1011
rect 730 1009 734 1010
rect 392 997 399 1001
rect 447 997 454 1001
rect 570 997 897 1001
rect 379 993 384 997
rect 380 987 384 989
rect 125 982 216 986
rect 125 973 129 982
rect 70 969 77 973
rect 125 969 132 973
rect -40 959 -36 968
rect -22 965 29 969
rect 34 965 62 969
rect -84 944 -58 949
rect -45 955 -36 959
rect 14 957 62 961
rect 70 957 74 969
rect 125 965 129 969
rect 117 961 129 965
rect -45 927 -40 955
rect 14 951 18 957
rect -159 926 -40 927
rect -220 925 -40 926
rect -214 922 -40 925
rect -31 947 18 951
rect -214 921 -154 922
rect -31 915 -27 947
rect 42 923 46 957
rect 70 953 77 957
rect 172 953 183 957
rect 65 949 74 953
rect 65 945 69 949
rect 212 948 216 982
rect 281 983 384 987
rect 392 985 396 997
rect 447 993 451 997
rect 439 989 451 993
rect 281 952 285 983
rect 392 981 399 985
rect 494 981 505 985
rect 387 977 396 981
rect 387 973 391 977
rect 226 948 233 952
rect 281 948 288 952
rect 212 944 218 948
rect 214 938 218 940
rect 132 936 218 938
rect 226 936 230 948
rect 281 944 285 948
rect 273 940 285 944
rect 132 934 217 936
rect 132 923 136 934
rect 42 919 136 923
rect -208 911 -27 915
rect -208 899 -204 911
rect -344 895 -204 899
rect 177 859 181 934
rect 226 932 233 936
rect 328 932 339 936
rect 221 928 230 932
rect 221 924 225 928
rect 570 874 574 997
rect 850 932 854 981
rect 905 941 909 1011
rect 941 1010 959 1011
rect 919 1002 959 1006
rect 967 1002 971 1014
rect 1022 1010 1026 1014
rect 1014 1006 1026 1010
rect 967 998 974 1002
rect 1069 998 1078 1002
rect 962 994 971 998
rect 962 991 966 994
rect 1821 984 1825 985
rect 1821 980 1923 984
rect 1821 974 1825 980
rect 1766 970 1773 974
rect 1821 970 1828 974
rect 1754 969 1758 970
rect 1598 966 1758 969
rect 1598 965 1757 966
rect 943 932 951 936
rect 994 932 1015 936
rect 595 927 615 931
rect 850 928 936 932
rect 597 921 601 927
rect 885 920 936 924
rect 943 920 948 932
rect 994 928 998 932
rect 991 924 998 928
rect 943 916 951 920
rect 910 912 936 916
rect 931 907 936 908
rect 605 874 609 881
rect 900 904 936 907
rect 943 904 948 916
rect 994 912 998 924
rect 1221 919 1497 923
rect 991 908 998 912
rect 900 903 935 904
rect 253 870 598 874
rect 605 870 847 874
rect 253 863 257 870
rect 605 867 609 870
rect 198 859 205 863
rect 253 859 260 863
rect 177 855 190 859
rect 189 847 190 851
rect 198 847 202 859
rect 253 855 257 859
rect 245 851 257 855
rect 198 843 205 847
rect 300 843 309 847
rect 671 865 675 870
rect 193 839 202 843
rect 597 843 601 847
rect 594 839 615 843
rect 193 836 197 839
rect 843 834 847 870
rect 900 820 904 903
rect 943 900 951 904
rect 943 890 948 900
rect 994 893 998 908
rect 1095 900 1116 904
rect 994 889 1150 893
rect 1146 883 1150 889
rect 1221 887 1225 919
rect 1493 897 1497 919
rect 1598 907 1602 965
rect 1665 958 1758 962
rect 1766 958 1770 970
rect 1821 966 1825 970
rect 1813 962 1825 966
rect 1665 922 1669 958
rect 1766 954 1773 958
rect 1868 954 1879 958
rect 1761 950 1770 954
rect 1761 946 1765 950
rect 1919 933 1923 980
rect 1987 937 1991 1030
rect 2170 1014 2174 1035
rect 2183 1027 2189 1032
rect 2185 1026 2189 1027
rect 2193 1026 2241 1029
rect 2212 1017 2216 1026
rect 2170 1010 2185 1014
rect 2181 1009 2185 1010
rect 1932 933 1939 937
rect 1987 933 1994 937
rect 1919 929 1924 933
rect 1920 923 1924 925
rect 1665 918 1756 922
rect 1665 909 1669 918
rect 1550 903 1602 907
rect 1610 905 1617 909
rect 1665 905 1672 909
rect 1598 901 1602 903
rect 1493 893 1602 897
rect 1610 893 1614 905
rect 1665 901 1669 905
rect 1657 897 1669 901
rect 1162 883 1170 887
rect 1213 883 1234 887
rect 1146 879 1155 883
rect 1010 871 1155 875
rect 1162 871 1167 883
rect 1213 879 1217 883
rect 1210 875 1217 879
rect 1010 839 1014 871
rect 1162 867 1170 871
rect 1130 863 1155 867
rect 1001 835 1019 839
rect 939 831 946 835
rect 954 827 961 831
rect 929 823 946 827
rect 556 819 942 820
rect 556 816 946 819
rect -147 773 -22 777
rect -456 769 -331 773
rect -456 761 -452 769
rect -513 757 -456 761
rect -537 752 -522 754
rect -547 750 -522 752
rect -547 748 -533 750
rect -513 736 -509 757
rect -500 749 -494 754
rect -498 748 -494 749
rect -490 748 -442 751
rect -471 737 -467 748
rect -513 732 -498 736
rect -502 731 -498 732
rect -446 724 -442 748
rect -446 719 -405 724
rect -456 710 -451 714
rect -456 705 -446 710
rect -450 704 -446 705
rect -417 668 -413 673
rect -438 664 -413 668
rect -486 635 -482 651
rect -467 652 -438 656
rect -467 635 -463 652
rect -494 631 -463 635
rect -494 615 -490 631
rect -417 609 -413 664
rect -410 657 -405 719
rect -399 708 -395 769
rect -337 767 -331 769
rect -337 763 -324 767
rect -387 719 -382 723
rect -399 704 -386 708
rect -337 698 -331 763
rect -147 765 -143 773
rect -204 761 -147 765
rect -228 756 -213 758
rect -238 754 -213 756
rect -238 752 -224 754
rect -204 740 -200 761
rect -191 753 -185 758
rect -189 752 -185 753
rect -181 752 -133 755
rect -162 741 -158 752
rect -204 736 -189 740
rect -193 735 -189 736
rect -337 694 -326 698
rect -330 690 -326 694
rect -382 660 -343 664
rect -410 656 -374 657
rect -410 652 -378 656
rect -450 599 -446 609
rect -434 605 -413 609
rect -347 642 -343 660
rect -137 728 -133 752
rect -137 723 -96 728
rect -147 714 -142 718
rect -147 709 -137 714
rect -141 708 -137 709
rect -108 672 -104 677
rect -129 668 -104 672
rect -337 642 -329 643
rect -502 592 -498 595
rect -450 594 -444 599
rect -504 587 -498 592
rect -504 577 -499 587
rect -510 574 -499 577
rect -449 575 -444 594
rect -390 575 -386 609
rect -374 597 -370 609
rect -353 639 -329 642
rect -322 642 -318 650
rect -353 637 -335 639
rect -322 638 -305 642
rect -177 639 -173 655
rect -158 656 -129 660
rect -158 639 -154 656
rect -353 597 -348 637
rect -322 636 -318 638
rect -330 607 -326 616
rect -374 592 -348 597
rect -335 603 -326 607
rect -335 575 -330 603
rect -449 574 -330 575
rect -510 573 -330 574
rect -504 570 -330 573
rect -504 569 -444 570
rect -309 551 -305 638
rect -185 635 -154 639
rect -185 619 -181 635
rect -108 613 -104 668
rect -101 661 -96 723
rect -90 712 -86 773
rect -28 771 -22 773
rect -28 767 -15 771
rect -78 723 -73 727
rect -90 708 -77 712
rect -28 702 -22 767
rect 556 728 560 816
rect 651 811 655 816
rect 843 755 847 808
rect 919 763 923 816
rect 938 815 946 816
rect 954 815 958 827
rect 1005 823 1009 835
rect 1001 819 1009 823
rect 954 811 961 815
rect 1079 811 1096 815
rect 954 805 958 811
rect 1130 788 1134 863
rect 1018 784 1134 788
rect 1146 855 1155 859
rect 1162 855 1167 867
rect 1213 863 1217 875
rect 1210 859 1217 863
rect 1018 766 1022 784
rect 919 762 949 763
rect 963 762 970 766
rect 1018 762 1025 766
rect 919 759 955 762
rect 945 758 955 759
rect 843 754 951 755
rect 843 751 955 754
rect 945 750 955 751
rect 963 750 967 762
rect 1018 758 1022 762
rect 1010 754 1022 758
rect 963 746 970 750
rect 1065 746 1074 750
rect 958 742 967 746
rect 958 739 962 742
rect 1146 738 1150 855
rect 1162 851 1170 855
rect 1314 851 1332 855
rect 1165 845 1169 851
rect 556 724 1123 728
rect 280 706 284 707
rect 280 702 382 706
rect -28 698 -17 702
rect -21 694 -17 698
rect 280 696 284 702
rect -73 664 -34 668
rect -101 660 -65 661
rect -101 656 -69 660
rect -141 603 -137 613
rect -125 609 -104 613
rect -38 646 -34 664
rect 225 692 232 696
rect 280 692 287 696
rect 213 691 217 692
rect -28 646 -20 647
rect -193 596 -189 599
rect -141 598 -135 603
rect -195 591 -189 596
rect -195 581 -190 591
rect -201 578 -190 581
rect -140 579 -135 598
rect -81 579 -77 613
rect -65 601 -61 613
rect -44 643 -20 646
rect -13 646 -9 654
rect 57 688 217 691
rect 57 687 216 688
rect -44 641 -26 643
rect -13 642 11 646
rect -44 601 -39 641
rect -13 640 -9 642
rect 7 627 11 642
rect 57 627 61 687
rect 124 680 217 684
rect 225 680 229 692
rect 280 688 284 692
rect 272 684 284 688
rect 124 644 128 680
rect 225 676 232 680
rect 327 676 338 680
rect 220 672 229 676
rect 220 668 224 672
rect 378 655 382 702
rect 556 673 560 724
rect 1144 721 1150 738
rect 1144 708 1148 721
rect 446 669 560 673
rect 590 704 1148 708
rect 446 659 450 669
rect 391 655 398 659
rect 446 655 453 659
rect 378 651 383 655
rect 379 645 383 647
rect 124 640 215 644
rect 124 631 128 640
rect 69 627 76 631
rect 124 627 131 631
rect 7 623 28 627
rect 33 623 61 627
rect -21 611 -17 620
rect -65 596 -39 601
rect -26 607 -17 611
rect 13 615 61 619
rect 69 615 73 627
rect 124 623 128 627
rect 116 619 128 623
rect 13 609 17 615
rect -26 579 -21 607
rect -140 578 -21 579
rect -201 577 -21 578
rect -195 574 -21 577
rect 7 605 17 609
rect -195 573 -135 574
rect 7 569 11 605
rect 41 581 45 615
rect 69 611 76 615
rect 171 611 182 615
rect 64 607 73 611
rect 64 603 68 607
rect 211 606 215 640
rect 280 641 383 645
rect 391 643 395 655
rect 446 651 450 655
rect 438 647 450 651
rect 590 648 594 704
rect 557 644 594 648
rect 280 610 284 641
rect 391 639 398 643
rect 493 639 504 643
rect 386 635 395 639
rect 386 631 390 635
rect 225 606 232 610
rect 280 606 287 610
rect 211 602 217 606
rect 213 596 217 598
rect 131 594 217 596
rect 225 594 229 606
rect 280 602 284 606
rect 272 598 284 602
rect 131 592 216 594
rect 131 581 135 592
rect 41 577 135 581
rect -191 565 11 569
rect -191 551 -187 565
rect -309 547 -187 551
rect 176 517 180 592
rect 225 590 232 594
rect 327 590 338 594
rect 220 586 229 590
rect 220 582 224 586
rect 557 532 561 644
rect 586 585 609 589
rect 591 579 595 585
rect 599 532 603 539
rect 252 528 592 532
rect 599 528 617 532
rect 252 521 256 528
rect 599 525 603 528
rect 197 517 204 521
rect 252 517 259 521
rect 176 513 189 517
rect 188 505 189 509
rect 197 505 201 517
rect 252 513 256 517
rect 244 509 256 513
rect 197 501 204 505
rect 299 501 308 505
rect 192 497 201 501
rect 591 501 595 505
rect 585 497 609 501
rect 192 494 196 497
rect -537 438 -412 442
rect -537 430 -533 438
rect -594 426 -537 430
rect -618 421 -603 423
rect -628 419 -603 421
rect -628 417 -614 419
rect -594 405 -590 426
rect -581 418 -575 423
rect -579 417 -575 418
rect -571 417 -523 420
rect -552 406 -548 417
rect -594 401 -579 405
rect -583 400 -579 401
rect -527 393 -523 417
rect -527 388 -486 393
rect -537 379 -532 383
rect -537 374 -527 379
rect -531 373 -527 374
rect -498 337 -494 342
rect -519 333 -494 337
rect -567 304 -563 320
rect -548 321 -519 325
rect -548 304 -544 321
rect -575 300 -544 304
rect -575 284 -571 300
rect -498 278 -494 333
rect -491 326 -486 388
rect -480 377 -476 438
rect -418 436 -412 438
rect -199 438 -74 442
rect -418 432 -405 436
rect -468 388 -463 392
rect -480 373 -467 377
rect -418 367 -412 432
rect -199 430 -195 438
rect -256 426 -199 430
rect -280 421 -265 423
rect -290 419 -265 421
rect -290 417 -276 419
rect -256 405 -252 426
rect -243 418 -237 423
rect -241 417 -237 418
rect -233 417 -185 420
rect -214 406 -210 417
rect -256 401 -241 405
rect -245 400 -241 401
rect -418 363 -407 367
rect -411 359 -407 363
rect -463 329 -424 333
rect -491 325 -455 326
rect -491 321 -459 325
rect -531 268 -527 278
rect -515 274 -494 278
rect -428 311 -424 329
rect -189 393 -185 417
rect -189 388 -148 393
rect -199 379 -194 383
rect -199 374 -189 379
rect -193 373 -189 374
rect -160 337 -156 342
rect -181 333 -156 337
rect -418 311 -410 312
rect -583 261 -579 264
rect -531 263 -525 268
rect -585 256 -579 261
rect -585 246 -580 256
rect -591 243 -580 246
rect -530 244 -525 263
rect -471 244 -467 278
rect -455 266 -451 278
rect -434 308 -410 311
rect -403 311 -399 319
rect -434 306 -416 308
rect -403 307 -369 311
rect -434 266 -429 306
rect -403 305 -399 307
rect -411 276 -407 285
rect -455 261 -429 266
rect -416 272 -407 276
rect -416 244 -411 272
rect -530 243 -411 244
rect -591 242 -411 243
rect -585 239 -411 242
rect -585 238 -525 239
rect -373 214 -369 307
rect -229 304 -225 320
rect -210 321 -181 325
rect -210 304 -206 321
rect -237 300 -206 304
rect -237 284 -233 300
rect -160 278 -156 333
rect -153 326 -148 388
rect -142 377 -138 438
rect -80 436 -74 438
rect -80 432 -67 436
rect -130 388 -125 392
rect -142 373 -129 377
rect -80 367 -74 432
rect 274 424 278 425
rect 274 420 376 424
rect 274 414 278 420
rect 219 410 226 414
rect 274 410 281 414
rect 207 409 211 410
rect 51 406 211 409
rect 51 405 210 406
rect -80 363 -69 367
rect -73 359 -69 363
rect -125 329 -86 333
rect -153 325 -117 326
rect -153 321 -121 325
rect -193 268 -189 278
rect -177 274 -156 278
rect -90 311 -86 329
rect 51 345 55 405
rect 118 398 211 402
rect 219 398 223 410
rect 274 406 278 410
rect 266 402 278 406
rect 118 362 122 398
rect 219 394 226 398
rect 321 394 332 398
rect 214 390 223 394
rect 214 386 218 390
rect 372 373 376 420
rect 613 404 617 528
rect 1545 524 1549 876
rect 1582 859 1586 893
rect 1610 889 1617 893
rect 1712 889 1723 893
rect 1605 885 1614 889
rect 1605 881 1609 885
rect 1752 884 1756 918
rect 1821 919 1924 923
rect 1932 921 1936 933
rect 1987 929 1991 933
rect 2237 1002 2241 1026
rect 2237 997 2278 1002
rect 2227 988 2232 992
rect 2227 983 2237 988
rect 2233 982 2237 983
rect 2266 946 2270 951
rect 2245 942 2270 946
rect 1979 925 1991 929
rect 1821 888 1825 919
rect 1932 917 1939 921
rect 2034 917 2045 921
rect 1927 913 1936 917
rect 2197 913 2201 929
rect 2216 930 2245 934
rect 2216 913 2220 930
rect 1927 909 1931 913
rect 2189 909 2220 913
rect 2189 893 2193 909
rect 1766 884 1773 888
rect 1821 884 1828 888
rect 1752 880 1758 884
rect 1754 874 1758 876
rect 1672 872 1758 874
rect 1766 872 1770 884
rect 1821 880 1825 884
rect 1813 876 1825 880
rect 2266 887 2270 942
rect 2273 935 2278 997
rect 2284 986 2288 1047
rect 2346 1043 2352 1047
rect 2346 1039 2359 1043
rect 2296 997 2301 1001
rect 2284 982 2297 986
rect 2346 976 2352 1039
rect 2346 972 2357 976
rect 2353 968 2357 972
rect 2301 938 2340 942
rect 2273 934 2309 935
rect 2273 930 2305 934
rect 2233 877 2237 887
rect 2249 883 2270 887
rect 2336 920 2340 938
rect 2346 920 2354 921
rect 1672 870 1757 872
rect 1672 859 1676 870
rect 1766 868 1773 872
rect 1868 868 1879 872
rect 2181 870 2185 873
rect 2233 872 2239 877
rect 1761 864 1770 868
rect 2179 865 2185 870
rect 1761 860 1765 864
rect 1582 855 1676 859
rect 2179 856 2184 865
rect 2173 852 2184 856
rect 2234 853 2239 872
rect 2293 853 2297 887
rect 2309 875 2313 887
rect 2330 917 2354 920
rect 2361 920 2365 928
rect 2330 915 2348 917
rect 2361 916 2371 920
rect 2330 875 2335 915
rect 2361 914 2365 916
rect 2353 885 2357 894
rect 2309 870 2335 875
rect 2348 881 2357 885
rect 2348 853 2353 881
rect 2234 852 2353 853
rect 2179 848 2353 852
rect 2179 847 2239 848
rect 632 520 1549 524
rect 632 391 636 520
rect 761 441 903 445
rect 899 426 903 441
rect 959 426 983 430
rect 899 422 904 426
rect 911 418 919 422
rect 815 414 904 418
rect 765 406 904 410
rect 911 406 915 418
rect 964 414 968 426
rect 959 410 968 414
rect 911 402 919 406
rect 664 398 904 402
rect 873 391 904 394
rect 440 390 904 391
rect 911 390 915 402
rect 964 398 968 410
rect 959 394 968 398
rect 440 387 877 390
rect 440 377 444 387
rect 385 373 392 377
rect 440 373 447 377
rect 550 376 554 387
rect 911 386 919 390
rect 911 377 915 386
rect 372 369 377 373
rect 373 363 377 365
rect 118 358 209 362
rect 118 349 122 358
rect 63 345 70 349
rect 118 345 125 349
rect -80 311 -72 312
rect -245 261 -241 264
rect -193 263 -187 268
rect -247 256 -241 261
rect -247 246 -242 256
rect -253 243 -242 246
rect -192 244 -187 263
rect -133 244 -129 278
rect -117 266 -113 278
rect -96 308 -72 311
rect -65 311 -61 319
rect -43 341 22 345
rect -43 311 -39 341
rect 27 341 55 345
rect 7 333 55 337
rect 63 333 67 345
rect 118 341 122 345
rect 110 337 122 341
rect 7 327 11 333
rect 1 323 11 327
rect -96 306 -78 308
rect -65 307 -39 311
rect -96 266 -91 306
rect -65 305 -61 307
rect -73 276 -69 285
rect -117 261 -91 266
rect -78 272 -69 276
rect -78 244 -73 272
rect -192 243 -73 244
rect -253 242 -73 243
rect -247 239 -73 242
rect -247 238 -187 239
rect 2 224 6 323
rect 35 299 39 333
rect 63 329 70 333
rect 165 329 176 333
rect 58 325 67 329
rect 58 321 62 325
rect 205 324 209 358
rect 274 359 377 363
rect 385 361 389 373
rect 440 369 444 373
rect 971 373 975 426
rect 1063 386 1083 390
rect 1670 386 1795 390
rect 1670 378 1674 386
rect 1613 374 1670 378
rect 971 369 1187 373
rect 1589 369 1604 371
rect 432 365 444 369
rect 274 328 278 359
rect 385 357 392 361
rect 487 357 498 361
rect 380 353 389 357
rect 380 349 384 353
rect 613 336 617 369
rect 1039 346 1166 350
rect 1162 333 1166 346
rect 1183 341 1187 369
rect 1256 367 1604 369
rect 1256 365 1593 367
rect 1256 345 1260 365
rect 1613 353 1617 374
rect 1626 366 1632 371
rect 1628 365 1632 366
rect 1636 365 1684 368
rect 1655 354 1659 365
rect 1613 349 1628 353
rect 1624 348 1628 349
rect 1243 341 1267 345
rect 1183 337 1188 341
rect 1195 333 1203 337
rect 1162 329 1188 333
rect 219 324 226 328
rect 274 324 281 328
rect 966 325 1136 329
rect 205 320 211 324
rect 207 314 211 316
rect 125 312 211 314
rect 219 312 223 324
rect 274 320 278 324
rect 266 316 278 320
rect 966 316 970 325
rect 1132 324 1136 325
rect 1183 324 1188 325
rect 1132 320 1188 324
rect 1195 321 1199 333
rect 1248 329 1252 341
rect 1243 325 1252 329
rect 1195 317 1203 321
rect 125 310 210 312
rect 125 299 129 310
rect 35 295 129 299
rect 170 235 174 310
rect 219 308 226 312
rect 321 308 332 312
rect 552 312 970 316
rect 1010 313 1188 317
rect 214 304 223 308
rect 214 300 218 304
rect 552 250 556 312
rect 993 305 1188 309
rect 1195 305 1199 317
rect 1248 313 1252 325
rect 1243 309 1252 313
rect 246 246 556 250
rect 246 239 250 246
rect 191 235 198 239
rect 246 235 253 239
rect 170 231 183 235
rect -236 220 6 224
rect 182 223 183 227
rect 191 223 195 235
rect 246 231 250 235
rect 238 227 250 231
rect -236 214 -232 220
rect 191 219 198 223
rect 293 219 302 223
rect -373 210 -232 214
rect 186 215 195 219
rect 186 212 190 215
rect 613 60 617 293
rect 703 268 925 272
rect 993 269 997 305
rect 1195 301 1203 305
rect 1347 301 1367 305
rect 1195 292 1199 301
rect 921 265 925 268
rect 933 265 941 269
rect 984 265 1005 269
rect 1680 341 1684 365
rect 1680 336 1721 341
rect 1670 327 1675 331
rect 1670 322 1680 327
rect 1676 321 1680 322
rect 1709 285 1713 290
rect 1688 281 1713 285
rect 921 261 926 265
rect 816 253 926 257
rect 933 253 938 265
rect 984 261 988 265
rect 981 257 988 261
rect 933 249 941 253
rect 857 245 926 249
rect 857 109 861 245
rect 905 237 926 241
rect 933 237 938 249
rect 984 245 988 257
rect 1640 252 1644 268
rect 1659 269 1688 273
rect 1659 252 1663 269
rect 1632 248 1663 252
rect 981 241 988 245
rect 905 106 909 237
rect 933 233 941 237
rect 1085 233 1103 237
rect 936 227 940 233
rect 1632 232 1636 248
rect 1709 226 1713 281
rect 1716 274 1721 336
rect 1727 325 1731 386
rect 1789 384 1795 386
rect 1789 380 1802 384
rect 1739 336 1744 340
rect 1727 321 1740 325
rect 1789 315 1795 380
rect 1789 311 1800 315
rect 1796 307 1800 311
rect 1744 277 1783 281
rect 1716 273 1752 274
rect 1716 269 1748 273
rect 1676 216 1680 226
rect 1692 222 1713 226
rect 1779 259 1783 277
rect 1789 259 1797 260
rect 1624 209 1628 212
rect 1676 211 1682 216
rect 1622 204 1628 209
rect 1622 194 1627 204
rect 1616 191 1627 194
rect 1677 192 1682 211
rect 1736 192 1740 226
rect 1752 214 1756 226
rect 1773 256 1797 259
rect 1804 259 1808 267
rect 1773 254 1791 256
rect 1804 255 1814 259
rect 1773 214 1778 254
rect 1804 253 1808 255
rect 1796 224 1800 233
rect 1752 209 1778 214
rect 1791 220 1800 224
rect 1791 192 1796 220
rect 1677 191 1796 192
rect 1616 190 1796 191
rect 1622 187 1796 190
rect 1622 186 1682 187
rect 1003 125 1007 139
rect 994 121 1012 125
rect 933 117 939 121
rect 947 113 954 117
rect 922 109 939 113
rect 905 105 935 106
rect 905 102 939 105
rect 613 56 873 60
rect 905 23 909 102
rect 932 101 939 102
rect 947 101 951 113
rect 998 109 1002 121
rect 994 105 1002 109
rect 947 97 954 101
rect 1072 97 1089 101
rect 947 91 951 97
rect 936 31 940 55
rect 1022 35 1026 50
rect 967 31 974 35
rect 1022 31 1029 35
rect 936 27 959 31
rect 895 19 959 23
rect 967 19 971 31
rect 1022 27 1026 31
rect 1014 23 1026 27
rect 967 15 974 19
rect 1069 15 1078 19
rect 962 11 971 15
rect 962 8 966 11
<< m2contact >>
rect -144 1882 -139 1887
rect -78 1889 -73 1894
rect -127 1882 -122 1887
rect -93 1865 -88 1870
rect -78 1847 -73 1852
rect -40 1806 -35 1811
rect -14 1852 -9 1857
rect 54 1895 59 1900
rect 658 1870 663 1875
rect -137 1705 -132 1710
rect 362 1710 367 1715
rect 243 1697 248 1702
rect 724 1877 729 1882
rect 675 1870 680 1875
rect 709 1856 714 1861
rect 724 1835 729 1840
rect 762 1794 767 1799
rect 788 1840 793 1845
rect 856 1883 861 1888
rect 665 1693 670 1698
rect 2156 1731 2161 1736
rect 52 1656 57 1661
rect -214 1632 -209 1637
rect -148 1639 -143 1644
rect -197 1632 -192 1637
rect -163 1615 -158 1620
rect -148 1597 -143 1602
rect -110 1556 -105 1561
rect -84 1602 -79 1607
rect -16 1645 -11 1650
rect -207 1455 -202 1460
rect 206 1645 211 1650
rect 87 1632 92 1637
rect 528 1673 533 1678
rect 409 1660 414 1665
rect 362 1624 367 1629
rect 606 1619 611 1624
rect 243 1611 248 1616
rect 1521 1576 1527 1582
rect 1870 1624 1875 1629
rect 1751 1611 1756 1616
rect 2222 1738 2227 1743
rect 2173 1731 2178 1736
rect 2204 1729 2210 1735
rect 2222 1696 2227 1701
rect 2260 1655 2265 1660
rect 207 1538 212 1543
rect 332 1535 337 1540
rect 604 1531 609 1536
rect 215 1523 220 1528
rect -539 1405 -534 1410
rect -473 1412 -468 1417
rect -522 1405 -517 1410
rect -488 1388 -483 1393
rect -473 1370 -468 1375
rect -435 1329 -430 1334
rect -409 1375 -404 1380
rect -341 1418 -336 1423
rect -182 1408 -177 1413
rect -116 1415 -111 1420
rect -165 1408 -160 1413
rect -131 1391 -126 1396
rect -116 1373 -111 1378
rect -78 1332 -73 1337
rect -532 1228 -527 1233
rect -52 1378 -47 1383
rect 16 1421 21 1426
rect 369 1359 374 1364
rect 250 1346 255 1351
rect 601 1352 606 1357
rect -175 1231 -170 1236
rect 59 1305 64 1310
rect 213 1294 218 1299
rect 94 1281 99 1286
rect 535 1322 540 1327
rect 416 1309 421 1314
rect 1714 1559 1719 1564
rect 1595 1546 1600 1551
rect 2036 1587 2041 1592
rect 1917 1574 1922 1579
rect 2286 1701 2291 1706
rect 2354 1747 2359 1752
rect 2163 1552 2168 1557
rect 1870 1538 1875 1543
rect 1751 1525 1756 1530
rect 2160 1471 2165 1476
rect 774 1310 779 1315
rect 923 1300 928 1305
rect 850 1285 855 1290
rect 932 1285 937 1290
rect 1075 1289 1080 1294
rect 369 1273 374 1278
rect 958 1277 963 1282
rect 609 1268 614 1273
rect 250 1260 255 1265
rect 1870 1349 1875 1354
rect 1751 1336 1756 1341
rect 2226 1478 2231 1483
rect 2177 1471 2182 1476
rect 2204 1469 2210 1475
rect 2226 1436 2231 1441
rect 2264 1395 2269 1400
rect 1535 1295 1540 1300
rect 1535 1269 1540 1274
rect 214 1187 219 1192
rect 339 1184 344 1189
rect 222 1172 227 1177
rect 862 1208 867 1213
rect 914 1211 919 1216
rect 684 1199 689 1204
rect 607 1180 612 1185
rect 651 1172 656 1177
rect 1001 1172 1006 1177
rect 1299 1224 1304 1229
rect 1182 1212 1187 1217
rect 651 1146 656 1151
rect 923 1149 928 1154
rect 932 1149 937 1154
rect 1001 1150 1006 1155
rect -563 1091 -558 1096
rect -497 1098 -492 1103
rect -546 1091 -541 1096
rect -512 1074 -507 1079
rect -497 1056 -492 1061
rect -459 1015 -454 1020
rect -433 1061 -428 1066
rect -365 1104 -360 1109
rect -232 1101 -227 1106
rect -166 1108 -161 1113
rect -215 1101 -210 1106
rect -181 1084 -176 1089
rect -166 1066 -161 1071
rect -128 1025 -123 1030
rect -556 914 -551 919
rect -102 1071 -97 1076
rect -34 1114 -29 1119
rect -225 924 -220 929
rect 339 1018 344 1023
rect 220 1005 225 1010
rect 1714 1284 1719 1289
rect 1595 1271 1600 1276
rect 2290 1441 2295 1446
rect 2358 1487 2363 1492
rect 2036 1312 2041 1317
rect 1917 1299 1922 1304
rect 2169 1295 2174 1300
rect 1870 1263 1875 1268
rect 1751 1250 1756 1255
rect 957 1063 962 1068
rect 1100 1074 1105 1079
rect 1554 1104 1559 1109
rect 1872 1155 1877 1160
rect 1753 1142 1758 1147
rect 2168 1247 2173 1252
rect 2234 1254 2239 1259
rect 2185 1247 2190 1252
rect 2214 1244 2220 1250
rect 2234 1212 2239 1217
rect 2272 1171 2277 1176
rect 1716 1090 1721 1095
rect 1597 1077 1602 1082
rect 2038 1118 2043 1123
rect 1919 1105 1924 1110
rect 2298 1217 2303 1222
rect 2366 1254 2371 1259
rect 1872 1069 1877 1074
rect 2175 1072 2180 1077
rect 1098 1037 1103 1042
rect 1753 1056 1758 1061
rect 1289 1033 1294 1038
rect 1146 1022 1151 1027
rect 725 1005 730 1010
rect 897 997 902 1002
rect 29 964 34 969
rect 183 953 188 958
rect 64 940 69 945
rect 505 981 510 986
rect 386 968 391 973
rect 339 932 344 937
rect 220 919 225 924
rect 850 981 855 986
rect 914 1002 919 1007
rect 1078 998 1083 1003
rect 961 986 966 991
rect 905 936 910 941
rect 590 927 595 932
rect 880 919 885 924
rect 905 911 910 916
rect 184 846 189 851
rect 309 843 314 848
rect 671 860 676 865
rect 589 839 594 844
rect 192 831 197 836
rect 843 829 848 834
rect 943 885 948 890
rect 1116 900 1121 905
rect 1879 954 1884 959
rect 1760 941 1765 946
rect 2161 1027 2166 1032
rect 2227 1034 2232 1039
rect 2178 1027 2183 1032
rect 2212 1012 2217 1017
rect 1545 902 1550 907
rect 1545 876 1550 881
rect 934 831 939 836
rect 924 823 929 828
rect -522 749 -517 754
rect -456 756 -451 761
rect -505 749 -500 754
rect -471 732 -466 737
rect -456 714 -451 719
rect -418 673 -413 678
rect -392 719 -387 724
rect -324 762 -319 767
rect -213 753 -208 758
rect -147 760 -142 765
rect -196 753 -191 758
rect -162 736 -157 741
rect -147 718 -142 723
rect -109 677 -104 682
rect -515 572 -510 577
rect -83 723 -78 728
rect -15 766 -10 771
rect 651 806 656 811
rect 843 808 848 813
rect 1096 811 1101 816
rect 953 800 958 805
rect 1074 746 1079 751
rect 957 734 962 739
rect 1332 851 1337 856
rect 1164 840 1169 845
rect 1123 724 1128 729
rect -206 576 -201 581
rect 338 676 343 681
rect 219 663 224 668
rect 28 622 33 627
rect 182 611 187 616
rect 63 598 68 603
rect 504 639 509 644
rect 385 626 390 631
rect 338 590 343 595
rect 219 577 224 582
rect 581 585 586 590
rect 183 504 188 509
rect 308 501 313 506
rect 580 497 585 502
rect 191 489 196 494
rect -603 418 -598 423
rect -537 425 -532 430
rect -586 418 -581 423
rect -552 401 -547 406
rect -537 383 -532 388
rect -499 342 -494 347
rect -473 388 -468 393
rect -405 431 -400 436
rect -265 418 -260 423
rect -199 425 -194 430
rect -248 418 -243 423
rect -214 401 -209 406
rect -199 383 -194 388
rect -161 342 -156 347
rect -596 241 -591 246
rect -135 388 -130 393
rect -67 431 -62 436
rect 332 394 337 399
rect 213 381 218 386
rect 1723 889 1728 894
rect 1604 876 1609 881
rect 2227 992 2232 997
rect 2265 951 2270 956
rect 2045 917 2050 922
rect 1926 904 1931 909
rect 2291 997 2296 1002
rect 2359 1038 2364 1043
rect 1879 868 1884 873
rect 1760 855 1765 860
rect 2168 851 2173 856
rect 613 399 618 404
rect 756 441 761 446
rect 815 418 820 423
rect 760 406 765 411
rect 659 398 664 403
rect -258 241 -253 246
rect 22 340 27 345
rect 176 329 181 334
rect 57 316 62 321
rect 550 371 555 376
rect 613 369 618 374
rect 910 372 915 377
rect 1083 386 1088 391
rect 498 357 503 362
rect 379 344 384 349
rect 1034 346 1039 351
rect 613 331 618 336
rect 1604 366 1609 371
rect 1670 373 1675 378
rect 1621 366 1626 371
rect 1655 349 1660 354
rect 332 308 337 313
rect 1005 312 1010 317
rect 213 295 218 300
rect 613 293 618 298
rect 177 222 182 227
rect 302 219 307 224
rect 185 207 190 212
rect 698 268 703 273
rect 1367 301 1372 306
rect 1194 287 1199 292
rect 1670 331 1675 336
rect 1708 290 1713 295
rect 811 253 816 259
rect 857 104 862 109
rect 1103 233 1108 238
rect 935 222 940 227
rect 1734 336 1739 341
rect 1802 379 1807 384
rect 1611 189 1616 194
rect 1003 139 1008 144
rect 928 117 933 122
rect 917 109 922 114
rect 873 56 878 61
rect 889 19 895 25
rect 1089 97 1094 102
rect 946 86 951 91
rect 936 55 941 60
rect 1022 50 1027 55
rect 1078 15 1083 20
rect 961 3 966 8
<< metal2 >>
rect 699 1941 2211 1945
rect 699 1923 703 1941
rect -174 1919 703 1923
rect -209 1632 -197 1636
rect -174 1609 -170 1919
rect -139 1882 -127 1886
rect -104 1859 -100 1919
rect 55 1890 59 1895
rect -93 1862 -88 1865
rect -93 1859 -82 1862
rect -104 1855 -82 1859
rect -101 1851 -82 1855
rect -78 1852 -73 1889
rect 663 1870 675 1874
rect -39 1852 -14 1856
rect -9 1852 -8 1856
rect -39 1811 -35 1852
rect 699 1851 703 1919
rect 857 1878 861 1883
rect 709 1851 713 1856
rect 699 1847 713 1851
rect 709 1846 713 1847
rect 724 1840 729 1877
rect 763 1840 788 1844
rect 793 1840 794 1844
rect 763 1799 767 1840
rect 2207 1830 2211 1941
rect 2205 1826 2211 1830
rect 2161 1731 2173 1735
rect 2205 1735 2209 1826
rect 2355 1742 2359 1747
rect 363 1715 367 1719
rect -137 1701 -133 1705
rect 238 1697 243 1701
rect 665 1689 669 1693
rect 529 1678 533 1682
rect 404 1660 409 1664
rect -15 1640 -11 1645
rect -163 1612 -158 1615
rect -163 1609 -152 1612
rect -174 1605 -152 1609
rect -171 1601 -152 1605
rect -148 1602 -143 1639
rect -207 1451 -203 1455
rect -162 1442 -158 1601
rect -109 1602 -84 1606
rect -79 1602 -78 1606
rect -109 1561 -105 1602
rect 52 1543 56 1656
rect 207 1650 211 1654
rect 82 1632 87 1636
rect 363 1629 367 1633
rect 1871 1629 1875 1633
rect 602 1619 606 1623
rect 238 1611 243 1615
rect 1746 1611 1751 1615
rect 2037 1592 2041 1596
rect 1327 1576 1521 1580
rect 52 1539 207 1543
rect 333 1540 337 1544
rect 600 1531 604 1535
rect 211 1523 215 1527
rect -142 1442 -138 1444
rect -499 1437 -263 1441
rect -534 1405 -522 1409
rect -499 1382 -495 1437
rect -267 1425 -263 1437
rect -191 1438 -138 1442
rect -191 1425 -187 1438
rect -267 1421 -187 1425
rect -340 1413 -336 1418
rect -488 1385 -483 1388
rect -488 1382 -477 1385
rect -499 1378 -477 1382
rect -496 1374 -477 1378
rect -473 1375 -468 1412
rect -177 1408 -165 1412
rect -142 1385 -138 1438
rect 17 1416 21 1421
rect -131 1388 -126 1391
rect -131 1385 -120 1388
rect -142 1381 -120 1385
rect -434 1375 -409 1379
rect -404 1375 -403 1379
rect -139 1377 -120 1381
rect -116 1378 -111 1415
rect -434 1334 -430 1375
rect -532 1224 -528 1228
rect -175 1227 -171 1231
rect -132 1169 -128 1377
rect -77 1378 -52 1382
rect -47 1378 -46 1382
rect -77 1337 -73 1378
rect 370 1364 374 1368
rect 1327 1356 1331 1576
rect 1912 1574 1917 1578
rect 1715 1564 1719 1568
rect 1590 1546 1595 1550
rect 1871 1543 1875 1547
rect 2163 1548 2167 1552
rect 1746 1525 1751 1529
rect 2165 1471 2177 1475
rect 2205 1475 2209 1729
rect 2222 1701 2227 1738
rect 2261 1701 2286 1705
rect 2291 1701 2292 1705
rect 2261 1660 2265 1701
rect 2359 1482 2363 1487
rect 606 1352 1331 1356
rect 1871 1354 1875 1358
rect 245 1346 250 1350
rect 1746 1336 1751 1340
rect 536 1327 540 1331
rect 746 1328 779 1332
rect 411 1309 416 1313
rect 59 1192 63 1305
rect 214 1299 218 1303
rect 89 1281 94 1285
rect 370 1278 374 1282
rect 605 1268 609 1272
rect 245 1260 250 1264
rect 59 1188 214 1192
rect 340 1189 344 1193
rect 603 1180 607 1184
rect 218 1172 222 1176
rect -234 1165 -128 1169
rect -234 1137 -230 1165
rect 651 1151 655 1172
rect -523 1133 -188 1137
rect -558 1091 -546 1095
rect -523 1068 -519 1133
rect -364 1099 -360 1104
rect -227 1101 -215 1105
rect -512 1071 -507 1074
rect -512 1068 -501 1071
rect -523 1064 -501 1068
rect -520 1060 -501 1064
rect -497 1061 -492 1098
rect -192 1078 -188 1133
rect -33 1109 -29 1114
rect -181 1081 -176 1084
rect -181 1078 -170 1081
rect -192 1074 -170 1078
rect -189 1070 -170 1074
rect -166 1071 -161 1108
rect -458 1061 -433 1065
rect -428 1061 -427 1065
rect -458 1020 -454 1061
rect -225 920 -221 924
rect -556 910 -552 914
rect -181 849 -177 1070
rect -127 1071 -102 1075
rect -97 1071 -96 1075
rect -127 1030 -123 1071
rect 340 1023 344 1027
rect 215 1005 220 1009
rect 506 986 510 990
rect -217 845 -177 849
rect 381 968 386 972
rect 29 851 33 964
rect 184 958 188 962
rect 59 940 64 944
rect 340 937 344 941
rect 586 927 590 931
rect 215 919 220 923
rect 29 847 184 851
rect 310 848 314 852
rect -217 801 -213 845
rect 585 839 589 843
rect 188 831 192 835
rect -483 797 -169 801
rect -483 785 -479 797
rect -483 777 -478 785
rect -517 749 -505 753
rect -482 726 -478 777
rect -323 757 -319 762
rect -471 729 -466 732
rect -471 726 -460 729
rect -482 722 -460 726
rect -479 718 -460 722
rect -456 719 -451 756
rect -208 753 -196 757
rect -173 730 -169 797
rect -14 761 -10 766
rect -162 733 -157 736
rect -162 730 -151 733
rect -173 726 -151 730
rect -417 719 -392 723
rect -387 719 -386 723
rect -170 722 -151 726
rect -147 723 -142 760
rect -417 678 -413 719
rect -206 572 -202 576
rect -515 568 -511 572
rect -164 488 -160 722
rect -108 723 -83 727
rect -78 723 -77 727
rect -108 682 -104 723
rect 339 681 343 685
rect 214 663 219 667
rect 505 644 509 648
rect 380 626 385 630
rect 28 509 32 622
rect 183 616 187 620
rect 58 598 63 602
rect 339 595 343 599
rect 577 585 581 589
rect 214 577 219 581
rect 28 505 183 509
rect 309 506 313 510
rect 576 497 580 501
rect 187 489 191 493
rect -239 484 -160 488
rect -239 462 -235 484
rect -563 458 -221 462
rect -598 418 -586 422
rect -563 395 -559 458
rect -404 426 -400 431
rect -552 398 -547 401
rect -552 395 -541 398
rect -563 391 -541 395
rect -560 387 -541 391
rect -537 388 -532 425
rect -260 418 -248 422
rect -225 395 -221 458
rect -66 426 -62 431
rect -214 398 -209 401
rect -214 395 -203 398
rect -498 388 -473 392
rect -468 388 -467 392
rect -225 391 -203 395
rect -498 347 -494 388
rect -222 387 -203 391
rect -199 388 -194 425
rect 333 399 337 403
rect 651 402 655 806
rect -160 388 -135 392
rect -130 388 -129 392
rect -160 347 -156 388
rect 208 381 213 385
rect 613 374 617 399
rect 651 398 659 402
rect 499 362 503 366
rect 374 344 379 348
rect -596 237 -592 241
rect -258 237 -254 241
rect 22 227 26 340
rect 177 334 181 338
rect 52 316 57 320
rect 333 313 337 317
rect 208 295 213 299
rect 22 223 177 227
rect 303 224 307 228
rect 181 207 185 211
rect 550 21 554 371
rect 613 298 617 331
rect 651 101 655 398
rect 671 124 675 860
rect 684 272 688 1199
rect 725 410 729 1005
rect 746 445 750 1328
rect 775 1315 779 1328
rect 2205 1325 2209 1469
rect 2226 1441 2231 1478
rect 2265 1441 2290 1445
rect 2295 1441 2296 1445
rect 2265 1400 2269 1441
rect 2205 1321 2219 1325
rect 2037 1317 2041 1321
rect 850 1075 854 1285
rect 923 1257 927 1300
rect 1076 1294 1080 1298
rect 880 1253 927 1257
rect 782 1071 854 1075
rect 746 441 756 445
rect 782 423 786 1071
rect 850 986 854 1071
rect 843 813 847 829
rect 862 827 866 1208
rect 880 924 884 1253
rect 914 1007 918 1211
rect 923 1154 927 1253
rect 1912 1299 1917 1303
rect 932 1154 936 1285
rect 954 1277 958 1281
rect 1535 1274 1539 1295
rect 1715 1289 1719 1293
rect 2169 1291 2173 1295
rect 1590 1271 1595 1275
rect 1871 1268 1875 1272
rect 1746 1250 1751 1254
rect 2173 1247 2185 1251
rect 2215 1250 2219 1321
rect 1300 1229 1304 1233
rect 1178 1212 1182 1216
rect 1001 1155 1005 1172
rect 1873 1160 1877 1164
rect 1748 1142 1753 1146
rect 2039 1123 2043 1127
rect 1388 1119 1542 1123
rect 1101 1079 1105 1083
rect 953 1063 957 1067
rect 923 1037 1098 1041
rect 1290 1038 1294 1042
rect 923 998 926 1037
rect 1142 1022 1146 1026
rect 1079 1003 1083 1007
rect 902 997 926 998
rect 897 994 926 997
rect 957 986 961 990
rect 905 916 909 936
rect 905 835 909 911
rect 1117 905 1121 909
rect 939 885 943 889
rect 1333 856 1337 860
rect 1160 840 1164 844
rect 905 832 934 835
rect 905 831 920 832
rect 933 831 934 832
rect 862 823 924 827
rect 1097 816 1101 820
rect 949 800 953 804
rect 1075 751 1079 755
rect 953 734 957 738
rect 1388 728 1392 1119
rect 1538 1108 1542 1119
rect 1538 1104 1554 1108
rect 1914 1105 1919 1109
rect 1717 1095 1721 1099
rect 2215 1085 2219 1244
rect 2234 1217 2239 1254
rect 2367 1249 2371 1254
rect 2273 1217 2298 1221
rect 2303 1217 2304 1221
rect 2273 1176 2277 1217
rect 1592 1077 1597 1081
rect 1873 1074 1877 1078
rect 2202 1081 2219 1085
rect 2175 1068 2179 1072
rect 1748 1056 1753 1060
rect 2166 1027 2178 1031
rect 2202 1010 2206 1081
rect 2211 1012 2212 1016
rect 2211 1010 2216 1012
rect 2202 1006 2216 1010
rect 1880 959 1884 963
rect 1755 941 1760 945
rect 2046 922 2050 926
rect 1921 904 1926 908
rect 1545 881 1549 902
rect 1724 894 1728 898
rect 1599 876 1604 880
rect 1880 873 1884 877
rect 1755 855 1760 859
rect 2168 847 2172 851
rect 2211 820 2215 1006
rect 2227 997 2232 1034
rect 2360 1033 2364 1038
rect 2266 997 2291 1001
rect 2296 997 2297 1001
rect 2266 956 2270 997
rect 1128 724 1392 728
rect 1644 816 2215 820
rect 782 419 815 423
rect 725 406 760 410
rect 684 268 698 272
rect 725 255 729 406
rect 1084 391 1088 395
rect 906 372 910 376
rect 1609 366 1621 370
rect 1022 346 1034 350
rect 1003 312 1005 317
rect 796 255 811 259
rect 725 251 800 255
rect 931 222 935 226
rect 1003 144 1007 312
rect 671 122 933 124
rect 671 120 928 122
rect 871 109 917 113
rect 871 105 875 109
rect 862 104 875 105
rect 857 101 875 104
rect 651 97 875 101
rect 942 86 946 90
rect 878 56 936 60
rect 1022 55 1026 346
rect 1644 343 1648 816
rect 1803 374 1807 379
rect 1655 346 1660 349
rect 1655 343 1666 346
rect 1644 339 1666 343
rect 1647 335 1666 339
rect 1670 336 1675 373
rect 1709 336 1734 340
rect 1739 336 1740 340
rect 1368 306 1372 310
rect 1709 295 1713 336
rect 1190 287 1194 291
rect 1104 238 1108 242
rect 1611 185 1615 189
rect 1090 102 1094 106
rect 550 19 889 21
rect 1079 20 1083 24
rect 550 17 893 19
rect 957 3 961 7
<< m3contact >>
rect 54 1885 59 1890
rect 856 1873 861 1878
rect 362 1719 367 1724
rect -137 1696 -132 1701
rect 233 1697 238 1702
rect 528 1682 533 1687
rect 665 1684 670 1689
rect 399 1660 404 1665
rect -16 1635 -11 1640
rect -207 1446 -202 1451
rect 206 1654 211 1659
rect 77 1632 82 1637
rect 362 1633 367 1638
rect 1870 1633 1875 1638
rect 597 1619 602 1624
rect 233 1611 238 1616
rect 1741 1611 1746 1616
rect 2036 1596 2041 1601
rect 332 1544 337 1549
rect 595 1531 600 1536
rect 206 1523 211 1528
rect -341 1408 -336 1413
rect 16 1411 21 1416
rect -532 1219 -527 1224
rect -175 1222 -170 1227
rect 369 1368 374 1373
rect 1907 1574 1912 1579
rect 1714 1568 1719 1573
rect 1585 1546 1590 1551
rect 1870 1547 1875 1552
rect 2163 1543 2168 1548
rect 1741 1525 1746 1530
rect 2354 1737 2359 1742
rect 1870 1358 1875 1363
rect 240 1346 245 1351
rect 1741 1336 1746 1341
rect 535 1331 540 1336
rect 406 1309 411 1314
rect 213 1303 218 1308
rect 84 1281 89 1286
rect 369 1282 374 1287
rect 600 1268 605 1273
rect 240 1260 245 1265
rect 339 1193 344 1198
rect 598 1180 603 1185
rect 213 1172 218 1177
rect -365 1094 -360 1099
rect -34 1104 -29 1109
rect -225 915 -220 920
rect -556 905 -551 910
rect 339 1027 344 1032
rect 210 1005 215 1010
rect 505 990 510 995
rect 376 968 381 973
rect 183 962 188 967
rect 54 940 59 945
rect 339 941 344 946
rect 581 927 586 932
rect 210 919 215 924
rect 309 852 314 857
rect 580 839 585 844
rect 183 831 188 836
rect -324 752 -319 757
rect -15 756 -10 761
rect -515 563 -510 568
rect -206 567 -201 572
rect 338 685 343 690
rect 209 663 214 668
rect 504 648 509 653
rect 375 626 380 631
rect 182 620 187 625
rect 53 598 58 603
rect 338 599 343 604
rect 572 585 577 590
rect 209 577 214 582
rect 308 510 313 515
rect 571 497 576 502
rect 182 489 187 494
rect -405 421 -400 426
rect -67 421 -62 426
rect 332 403 337 408
rect 203 381 208 386
rect 498 366 503 371
rect 369 344 374 349
rect -596 232 -591 237
rect -258 232 -253 237
rect 176 338 181 343
rect 47 316 52 321
rect 332 317 337 322
rect 203 295 208 300
rect 302 228 307 233
rect 176 207 181 212
rect 2036 1321 2041 1326
rect 2358 1477 2363 1482
rect 1075 1298 1080 1303
rect 1907 1299 1912 1304
rect 949 1277 954 1282
rect 1714 1293 1719 1298
rect 2169 1286 2174 1291
rect 1585 1271 1590 1276
rect 1870 1272 1875 1277
rect 1741 1250 1746 1255
rect 1299 1233 1304 1238
rect 1173 1212 1178 1217
rect 1872 1164 1877 1169
rect 1743 1142 1748 1147
rect 2038 1127 2043 1132
rect 1100 1083 1105 1088
rect 948 1063 953 1068
rect 1289 1042 1294 1047
rect 1137 1022 1142 1027
rect 1078 1007 1083 1012
rect 952 986 957 991
rect 1116 909 1121 914
rect 934 885 939 890
rect 1332 860 1337 865
rect 1155 840 1160 845
rect 1096 820 1101 825
rect 944 800 949 805
rect 1074 755 1079 760
rect 948 734 953 739
rect 1909 1105 1914 1110
rect 1716 1099 1721 1104
rect 2366 1244 2371 1249
rect 1587 1077 1592 1082
rect 1872 1078 1877 1083
rect 2175 1063 2180 1068
rect 1743 1056 1748 1061
rect 1879 963 1884 968
rect 1750 941 1755 946
rect 2045 926 2050 931
rect 1916 904 1921 909
rect 1723 898 1728 903
rect 1594 876 1599 881
rect 1879 877 1884 882
rect 1750 855 1755 860
rect 2168 842 2173 847
rect 2359 1028 2364 1033
rect 1083 395 1088 400
rect 901 372 906 377
rect 926 222 931 227
rect 937 86 942 91
rect 1802 369 1807 374
rect 1367 310 1372 315
rect 1185 287 1190 292
rect 1103 242 1108 247
rect 1611 180 1616 185
rect 1089 106 1094 111
rect 1078 24 1083 29
rect 952 3 957 8
<< metal3 >>
rect 36 1918 98 1922
rect 36 1887 40 1918
rect 36 1885 54 1887
rect 36 1883 59 1885
rect 94 1743 98 1918
rect 838 1918 892 1922
rect 838 1875 842 1918
rect 838 1873 856 1875
rect 838 1871 861 1873
rect 75 1742 235 1743
rect 75 1739 401 1742
rect -137 1692 -133 1696
rect 75 1672 79 1739
rect -34 1668 79 1672
rect -34 1637 -30 1668
rect -34 1635 -16 1637
rect -34 1633 -11 1635
rect 75 1637 79 1668
rect 75 1632 77 1637
rect 112 1458 116 1739
rect 172 1597 176 1739
rect 231 1738 401 1739
rect 231 1702 235 1738
rect 363 1724 367 1728
rect 231 1697 233 1702
rect 397 1667 401 1738
rect 529 1687 533 1691
rect 665 1680 669 1684
rect 397 1665 402 1667
rect 397 1664 399 1665
rect 207 1659 211 1663
rect 231 1660 399 1664
rect 231 1619 235 1660
rect 363 1638 367 1642
rect 554 1619 597 1623
rect 231 1616 236 1619
rect 231 1611 233 1616
rect 554 1597 558 1619
rect 172 1593 558 1597
rect 172 1532 176 1593
rect 333 1549 337 1553
rect 172 1528 210 1532
rect 587 1531 595 1535
rect 887 1458 891 1918
rect 1893 1776 2325 1780
rect 1583 1656 1743 1657
rect 1893 1656 1897 1776
rect 2321 1739 2325 1776
rect 2321 1737 2354 1739
rect 2321 1735 2359 1737
rect 1583 1653 1909 1656
rect 1583 1551 1587 1653
rect 1583 1546 1585 1551
rect 112 1454 1130 1458
rect -207 1442 -203 1446
rect -2 1443 2 1444
rect 112 1443 116 1454
rect -359 1431 -355 1441
rect -2 1439 116 1443
rect -2 1431 2 1439
rect -359 1427 2 1431
rect -359 1410 -355 1427
rect -2 1413 2 1427
rect -359 1408 -341 1410
rect -2 1411 16 1413
rect -2 1409 21 1411
rect -359 1406 -336 1408
rect 112 1392 116 1439
rect 1126 1448 1130 1454
rect 1625 1448 1629 1653
rect 1739 1652 1909 1653
rect 1739 1616 1743 1652
rect 1871 1638 1875 1642
rect 1739 1611 1741 1616
rect 1905 1581 1909 1652
rect 2037 1601 2041 1605
rect 1905 1579 1910 1581
rect 1905 1578 1907 1579
rect 1715 1573 1719 1577
rect 1739 1574 1907 1578
rect 1739 1533 1743 1574
rect 1871 1552 1875 1556
rect 2163 1539 2167 1543
rect 1739 1530 1744 1533
rect 1739 1525 1741 1530
rect 2325 1479 2329 1735
rect 2325 1477 2358 1479
rect 2325 1475 2363 1477
rect 1126 1444 1629 1448
rect 82 1391 242 1392
rect 82 1388 408 1391
rect 82 1286 86 1388
rect 82 1281 84 1286
rect -532 1215 -528 1219
rect -175 1218 -171 1222
rect -52 1128 -48 1137
rect 112 1128 116 1388
rect 179 1181 183 1388
rect 238 1387 408 1388
rect 238 1351 242 1387
rect 370 1373 374 1377
rect 238 1346 240 1351
rect 404 1316 408 1387
rect 536 1336 540 1340
rect 404 1314 409 1316
rect 404 1313 406 1314
rect 214 1308 218 1312
rect 238 1309 406 1313
rect 238 1273 242 1309
rect 1076 1303 1080 1307
rect 370 1287 374 1291
rect 941 1282 953 1286
rect 238 1272 253 1273
rect 238 1269 600 1272
rect 238 1265 243 1269
rect 249 1268 600 1269
rect 238 1260 240 1265
rect 941 1222 945 1282
rect 1126 1222 1130 1444
rect 1625 1382 1629 1444
rect 1583 1381 1743 1382
rect 1583 1378 1909 1381
rect 1583 1276 1587 1378
rect 1583 1271 1585 1276
rect 1300 1238 1304 1242
rect 941 1218 1178 1222
rect 340 1198 344 1202
rect 179 1177 217 1181
rect 590 1180 598 1184
rect -383 1123 116 1128
rect -383 1096 -379 1123
rect -52 1106 -48 1123
rect -52 1104 -34 1106
rect -52 1102 -29 1104
rect -383 1094 -365 1096
rect -383 1092 -360 1094
rect 112 1051 116 1123
rect 944 1073 948 1218
rect 1101 1088 1105 1092
rect 944 1068 952 1073
rect 52 1050 212 1051
rect 52 1047 378 1050
rect 52 945 56 1047
rect 52 940 54 945
rect -225 911 -221 915
rect -556 901 -552 905
rect -342 784 -338 785
rect -33 784 -29 789
rect 112 784 116 1047
rect 149 899 153 1047
rect 208 1046 378 1047
rect 208 1010 212 1046
rect 340 1032 344 1036
rect 208 1005 210 1010
rect 374 975 378 1046
rect 944 1033 948 1068
rect 1137 1033 1141 1218
rect 1164 1217 1178 1218
rect 1164 1216 1173 1217
rect 1625 1188 1629 1378
rect 1739 1377 1909 1378
rect 1739 1341 1743 1377
rect 1871 1363 1875 1367
rect 1739 1336 1741 1341
rect 1905 1306 1909 1377
rect 2037 1326 2041 1330
rect 1905 1304 1910 1306
rect 1905 1303 1907 1304
rect 1715 1298 1719 1302
rect 1739 1299 1907 1303
rect 1739 1258 1743 1299
rect 1871 1277 1875 1281
rect 2169 1282 2173 1286
rect 1739 1255 1744 1258
rect 1739 1250 1741 1255
rect 2338 1246 2342 1475
rect 2338 1244 2366 1246
rect 2338 1242 2371 1244
rect 1585 1187 1745 1188
rect 1585 1184 1911 1187
rect 1585 1082 1589 1184
rect 1585 1077 1587 1082
rect 1290 1047 1294 1051
rect 944 1029 1141 1033
rect 506 995 510 999
rect 944 995 948 1029
rect 1137 1027 1141 1029
rect 1079 1012 1083 1016
rect 1137 1016 1141 1022
rect 1137 1012 1159 1016
rect 944 994 957 995
rect 926 991 957 994
rect 926 990 952 991
rect 374 973 379 975
rect 374 972 376 973
rect 184 967 188 971
rect 208 968 376 972
rect 208 927 212 968
rect 340 946 344 950
rect 522 927 581 931
rect 208 924 213 927
rect 208 919 210 924
rect 522 899 526 927
rect 148 895 526 899
rect 149 840 153 895
rect 926 894 930 990
rect 1117 914 1121 918
rect 926 890 939 894
rect 933 889 934 890
rect 934 881 938 885
rect 934 877 944 881
rect 310 857 314 861
rect 149 836 187 840
rect 572 839 580 843
rect 940 810 944 877
rect 1155 845 1159 1012
rect 1625 987 1629 1184
rect 1741 1183 1911 1184
rect 1741 1147 1745 1183
rect 1873 1169 1877 1173
rect 1741 1142 1743 1147
rect 1907 1112 1911 1183
rect 2039 1132 2043 1136
rect 1907 1110 1912 1112
rect 1907 1109 1909 1110
rect 1717 1104 1721 1108
rect 1741 1105 1909 1109
rect 1741 1064 1745 1105
rect 1873 1083 1877 1087
rect 1741 1061 1746 1064
rect 1741 1056 1743 1061
rect 2175 1059 2179 1063
rect 2338 1030 2342 1242
rect 2338 1028 2359 1030
rect 2338 1026 2364 1028
rect 1592 986 1752 987
rect 1592 983 1918 986
rect 1592 881 1596 983
rect 1748 982 1918 983
rect 1748 946 1752 982
rect 1880 968 1884 972
rect 1748 941 1750 946
rect 1914 911 1918 982
rect 2046 931 2050 935
rect 1914 909 1919 911
rect 1914 908 1916 909
rect 1724 903 1728 907
rect 1748 904 1916 908
rect 1592 876 1594 881
rect 1333 865 1337 869
rect 1748 863 1752 904
rect 1880 882 1884 886
rect 1748 860 1753 863
rect 1748 855 1750 860
rect 2168 838 2172 842
rect 1097 825 1101 829
rect 940 805 948 810
rect 940 800 944 805
rect -342 780 116 784
rect -342 754 -338 780
rect -33 758 -29 780
rect -342 752 -324 754
rect -33 756 -15 758
rect -33 754 -10 756
rect -342 750 -319 752
rect 112 709 116 780
rect 945 775 949 800
rect 943 743 949 775
rect 1075 760 1079 764
rect 943 739 953 743
rect 943 734 948 739
rect 943 731 951 734
rect 51 708 211 709
rect 51 705 377 708
rect 51 603 55 705
rect 51 598 53 603
rect -206 563 -202 567
rect -515 559 -511 563
rect 112 454 116 705
rect 148 564 152 705
rect 207 704 377 705
rect 207 668 211 704
rect 339 690 343 694
rect 207 663 209 668
rect 373 633 377 704
rect 943 677 947 731
rect 882 673 947 677
rect 505 653 509 657
rect 373 631 378 633
rect 373 630 375 631
rect 183 625 187 629
rect 207 626 375 630
rect 207 585 211 626
rect 339 604 343 608
rect 549 585 572 589
rect 207 582 212 585
rect 207 577 209 582
rect 549 564 553 585
rect 148 560 553 564
rect 148 498 152 560
rect 309 515 313 519
rect 148 494 186 498
rect 563 497 571 501
rect -423 450 116 454
rect -423 423 -419 450
rect -423 421 -405 423
rect -423 419 -400 421
rect -85 423 -81 450
rect 112 427 116 450
rect 45 426 205 427
rect -85 421 -67 423
rect -85 419 -62 421
rect 45 423 371 426
rect 45 321 49 423
rect 45 316 47 321
rect -596 228 -592 232
rect -258 228 -254 232
rect 142 216 146 423
rect 201 422 371 423
rect 201 386 205 422
rect 333 408 337 412
rect 201 381 203 386
rect 367 351 371 422
rect 882 385 886 673
rect 1784 414 1878 418
rect 1084 400 1088 404
rect 882 381 902 385
rect 499 371 503 375
rect 367 349 372 351
rect 367 348 369 349
rect 177 343 181 347
rect 201 344 369 348
rect 201 303 205 344
rect 333 322 337 326
rect 201 300 206 303
rect 201 295 203 300
rect 882 296 886 381
rect 898 377 906 381
rect 898 376 901 377
rect 1784 371 1788 414
rect 1784 369 1802 371
rect 1784 367 1807 369
rect 1368 315 1372 319
rect 1182 296 1186 300
rect 882 292 1190 296
rect 303 233 307 237
rect 142 212 180 216
rect 902 207 906 292
rect 926 227 930 292
rect 1104 247 1108 251
rect 902 203 937 207
rect 933 96 937 203
rect 1149 126 1153 292
rect 1182 291 1185 292
rect 1611 176 1615 180
rect 1874 126 1878 414
rect 1149 122 1878 126
rect 1090 111 1094 115
rect 933 95 941 96
rect 922 91 941 95
rect 922 13 926 91
rect 933 86 937 91
rect 938 85 942 86
rect 1079 29 1083 33
rect 922 9 957 13
rect 943 8 957 9
rect 943 7 952 8
<< m4contact >>
rect -137 1687 -132 1692
rect 362 1728 367 1733
rect 206 1663 211 1668
rect 528 1691 533 1696
rect 665 1675 670 1680
rect 362 1642 367 1647
rect 332 1553 337 1558
rect 582 1530 587 1535
rect -207 1437 -202 1442
rect 1870 1642 1875 1647
rect 1714 1577 1719 1582
rect 2036 1605 2041 1610
rect 1870 1556 1875 1561
rect 2163 1534 2168 1539
rect -532 1210 -527 1215
rect -175 1213 -170 1218
rect 369 1377 374 1382
rect 213 1312 218 1317
rect 535 1340 540 1345
rect 1075 1307 1080 1312
rect 369 1291 374 1296
rect 1299 1242 1304 1247
rect 339 1202 344 1207
rect 585 1179 590 1184
rect 1100 1092 1105 1097
rect -225 906 -220 911
rect -556 896 -551 901
rect 339 1036 344 1041
rect 183 971 188 976
rect 1870 1367 1875 1372
rect 1714 1302 1719 1307
rect 2036 1330 2041 1335
rect 1870 1281 1875 1286
rect 2169 1277 2174 1282
rect 1289 1051 1294 1056
rect 505 999 510 1004
rect 1078 1016 1083 1021
rect 339 950 344 955
rect 1116 918 1121 923
rect 309 861 314 866
rect 567 838 572 843
rect 1872 1173 1877 1178
rect 1716 1108 1721 1113
rect 2038 1136 2043 1141
rect 1872 1087 1877 1092
rect 2175 1054 2180 1059
rect 1879 972 1884 977
rect 1723 907 1728 912
rect 2045 935 2050 940
rect 1332 869 1337 874
rect 1879 886 1884 891
rect 1096 829 1101 834
rect 2168 833 2173 838
rect 1074 764 1079 769
rect -515 554 -510 559
rect -206 558 -201 563
rect 338 694 343 699
rect 182 629 187 634
rect 504 657 509 662
rect 338 608 343 613
rect 308 519 313 524
rect 558 496 563 501
rect -596 223 -591 228
rect -258 223 -253 228
rect 332 412 337 417
rect 176 347 181 352
rect 1083 404 1088 409
rect 498 375 503 380
rect 332 326 337 331
rect 1367 319 1372 324
rect 302 237 307 242
rect 1103 251 1108 256
rect 1611 171 1616 176
rect 1089 115 1094 120
rect 1078 33 1083 38
<< metal4 >>
rect 367 1729 375 1733
rect -246 1687 -137 1691
rect -246 1584 -242 1687
rect 371 1668 375 1729
rect 533 1692 541 1696
rect 211 1664 375 1668
rect 371 1647 375 1664
rect 367 1646 375 1647
rect 537 1679 541 1692
rect 537 1675 665 1679
rect 537 1646 541 1675
rect 367 1643 541 1646
rect 371 1642 541 1643
rect 1875 1643 1883 1647
rect 384 1584 388 1642
rect -246 1580 388 1584
rect -246 1441 -242 1580
rect 384 1558 388 1580
rect 337 1554 388 1558
rect 448 1533 452 1642
rect 1879 1582 1883 1643
rect 2041 1606 2049 1610
rect 1719 1578 1883 1582
rect 1879 1561 1883 1578
rect 1875 1560 1883 1561
rect 2045 1560 2049 1606
rect 1875 1557 2049 1560
rect 1879 1556 2049 1557
rect 1979 1538 1983 1556
rect 580 1533 582 1535
rect 448 1530 582 1533
rect 1979 1534 2163 1538
rect 448 1529 584 1530
rect -246 1437 -207 1441
rect -246 1217 -242 1437
rect 448 1423 452 1529
rect 448 1419 1180 1423
rect 374 1378 382 1382
rect 378 1317 382 1378
rect 218 1313 382 1317
rect 378 1296 382 1313
rect 374 1295 382 1296
rect 448 1295 452 1419
rect 1176 1411 1180 1419
rect 1979 1411 1983 1534
rect 1176 1407 1983 1411
rect 540 1341 548 1345
rect 544 1295 548 1341
rect 1176 1312 1180 1407
rect 1875 1368 1883 1372
rect 1080 1308 1311 1312
rect 374 1292 548 1295
rect 378 1291 548 1292
rect -564 1210 -532 1214
rect -511 1213 -175 1217
rect -564 1203 -560 1210
rect -511 1203 -507 1213
rect -564 1199 -507 1203
rect -319 909 -315 1213
rect 391 1207 395 1291
rect 344 1203 395 1207
rect 448 1184 452 1291
rect 448 1179 585 1184
rect 344 1037 352 1041
rect 348 976 352 1037
rect 188 972 352 976
rect 348 955 352 972
rect 344 954 352 955
rect 448 954 452 1179
rect 1108 1097 1112 1308
rect 1307 1247 1311 1308
rect 1879 1307 1883 1368
rect 1719 1303 1883 1307
rect 1879 1286 1883 1303
rect 1875 1285 1883 1286
rect 1979 1285 1983 1407
rect 2041 1331 2049 1335
rect 2045 1285 2049 1331
rect 1875 1282 2049 1285
rect 1879 1281 2049 1282
rect 1304 1243 1311 1247
rect 1308 1239 1344 1243
rect 1105 1094 1113 1097
rect 1105 1093 1301 1094
rect 1109 1090 1301 1093
rect 1121 1021 1125 1090
rect 1297 1056 1301 1090
rect 1294 1052 1301 1056
rect 1083 1017 1128 1021
rect 510 1000 518 1004
rect 514 954 518 1000
rect 344 951 518 954
rect 348 950 518 951
rect -257 909 -225 910
rect -527 906 -225 909
rect -527 905 -252 906
rect -588 896 -556 900
rect -588 885 -584 896
rect -527 885 -523 905
rect -588 881 -523 885
rect -288 561 -284 905
rect 361 866 365 950
rect 314 862 365 866
rect 448 843 452 950
rect 1124 923 1128 1017
rect 1121 919 1128 923
rect 1125 914 1128 919
rect 448 839 567 843
rect 343 695 351 699
rect 347 634 351 695
rect 187 630 351 634
rect 347 613 351 630
rect 343 612 351 613
rect 448 612 452 839
rect 1124 834 1128 914
rect 1340 874 1344 1239
rect 1877 1174 1885 1178
rect 1881 1113 1885 1174
rect 1721 1109 1885 1113
rect 1881 1092 1885 1109
rect 1877 1091 1885 1092
rect 1979 1091 1983 1281
rect 2045 1277 2169 1281
rect 2043 1137 2051 1141
rect 2047 1091 2051 1137
rect 1877 1088 2051 1091
rect 1881 1087 2051 1088
rect 1979 1058 1983 1087
rect 1979 1054 2175 1058
rect 1884 973 1892 977
rect 1888 912 1892 973
rect 1728 908 1892 912
rect 1888 891 1892 908
rect 1884 890 1892 891
rect 1979 890 1983 1054
rect 2050 936 2058 940
rect 2054 890 2058 936
rect 1884 887 2058 890
rect 1888 886 2058 887
rect 1337 870 1344 874
rect 1101 830 1128 834
rect 2050 837 2054 886
rect 2050 833 2168 837
rect 1119 769 1123 830
rect 1079 767 1123 769
rect 1079 765 1303 767
rect 1117 763 1303 765
rect 509 658 517 662
rect 513 612 517 658
rect 343 609 517 612
rect 347 608 517 609
rect -238 561 -206 562
rect -547 554 -515 558
rect -496 558 -206 561
rect -496 557 -233 558
rect -547 544 -543 554
rect -496 544 -492 557
rect -547 540 -492 544
rect -628 223 -596 227
rect -288 227 -284 557
rect 360 524 364 608
rect 313 520 364 524
rect 448 501 452 608
rect 448 497 558 501
rect 337 413 345 417
rect 341 352 345 413
rect 181 348 345 352
rect 341 331 345 348
rect 337 330 345 331
rect 448 330 452 497
rect 1299 409 1303 763
rect 1088 405 1395 409
rect 503 376 511 380
rect 507 330 511 376
rect 337 327 511 330
rect 341 326 511 327
rect 354 242 358 326
rect 1111 265 1115 405
rect 1372 323 1376 324
rect 1391 323 1395 405
rect 1372 320 1395 323
rect 1380 319 1395 320
rect 1111 261 1129 265
rect 1111 256 1115 261
rect 1108 252 1115 256
rect 307 238 358 242
rect -573 223 -258 227
rect -625 213 -621 223
rect -573 213 -569 223
rect 1125 220 1129 261
rect -625 209 -569 213
rect 1096 216 1129 220
rect 1096 175 1100 216
rect 1096 171 1611 175
rect 1096 126 1100 171
rect 1096 122 1113 126
rect 1096 120 1100 122
rect 1094 116 1100 120
rect 1109 51 1113 122
rect 1086 47 1113 51
rect 1086 38 1090 47
rect 1083 34 1090 38
<< labels >>
rlabel metal1 582 1562 586 1566 1 gn0
rlabel metal1 587 1352 591 1356 7 p1
rlabel metal1 589 1211 593 1215 7 gn1
rlabel metal1 557 1011 561 1015 1 p2
rlabel metal1 559 870 563 874 1 gn2
rlabel metal1 556 669 560 673 1 p3
rlabel metal1 558 528 562 532 1 gn3
rlabel metal1 550 387 554 391 1 p4
rlabel metal1 552 246 556 250 1 gn4
rlabel metal1 637 1562 641 1566 7 g0
rlabel metal1 640 1211 644 1215 7 g1
rlabel metal1 619 870 623 874 1 g2
rlabel metal1 613 528 617 532 1 g3
rlabel metal1 1493 919 1497 923 1 c4
rlabel metal1 1489 1105 1493 1109 1 c3
rlabel metal1 1487 1264 1491 1268 1 c2
rlabel metal1 1480 1561 1484 1565 1 c1
rlabel metal3 146 1739 150 1743 5 vdd
rlabel metal4 537 1655 541 1659 1 gnd
rlabel metal1 2362 1620 2366 1624 1 s1
rlabel metal1 2366 1360 2370 1364 1 s2
rlabel metal1 2374 1136 2378 1140 7 s3
rlabel metal1 2367 916 2371 920 1 s4
rlabel metal1 1810 255 1814 259 1 cout
rlabel metal1 864 1759 868 1763 1 s0
rlabel metal2 1032 1941 1036 1945 5 clk
rlabel metal1 -152 1883 -148 1887 1 a0
rlabel metal1 -221 1633 -217 1637 1 b0
rlabel metal1 -207 1407 -203 1411 1 a1
rlabel metal1 -564 1404 -560 1408 1 b1
rlabel metal1 -257 1100 -253 1104 1 a2
rlabel metal1 -588 1090 -584 1094 1 b2
rlabel metal1 -238 752 -234 756 1 a3
rlabel metal1 -547 748 -543 752 1 b3
rlabel metal1 -276 419 -272 423 1 a4
rlabel metal1 -628 417 -624 421 3 b4
<< end >>
