magic
tech scmos
timestamp 1763472339
<< nwell >>
rect 147 978 199 1010
rect -9 913 43 945
rect 313 941 365 973
rect 147 892 199 924
rect 506 841 530 897
rect 1655 892 1707 924
rect 119 803 171 835
rect 1499 827 1551 859
rect 1821 855 1873 887
rect 1655 806 1707 838
rect 154 627 206 659
rect -2 562 50 594
rect 320 590 372 622
rect 1655 617 1707 649
rect 154 541 206 573
rect 862 557 914 589
rect 1499 552 1551 584
rect 1821 580 1873 612
rect 509 490 533 546
rect 1655 531 1707 563
rect 1086 492 1138 524
rect 126 452 178 484
rect 1657 423 1709 455
rect 856 354 908 382
rect 1501 358 1553 390
rect 1823 386 1875 418
rect 855 342 908 354
rect 124 286 176 318
rect 1045 313 1097 341
rect 1657 337 1709 369
rect 1044 301 1097 313
rect -32 221 20 253
rect 290 249 342 281
rect 865 266 917 298
rect 124 200 176 232
rect 1664 222 1716 254
rect 488 149 512 205
rect 842 168 894 216
rect 96 111 148 143
rect 1061 119 1113 167
rect 1508 157 1560 189
rect 1830 185 1882 217
rect 1664 136 1716 168
rect 852 91 904 119
rect 851 79 904 91
rect 861 14 913 46
rect 123 -56 175 -24
rect -33 -121 19 -89
rect 289 -93 341 -61
rect 123 -142 175 -110
rect 482 -193 506 -137
rect 95 -231 147 -199
rect 117 -338 169 -306
rect -39 -403 13 -371
rect 283 -375 335 -343
rect 810 -346 862 -290
rect 117 -424 169 -392
rect 1094 -431 1146 -375
rect 89 -513 141 -481
rect 832 -499 884 -451
rect 845 -623 897 -595
rect 844 -635 897 -623
rect 865 -717 917 -685
<< ntransistor >>
rect 208 997 248 999
rect 208 989 248 991
rect 374 960 414 962
rect 374 952 414 954
rect 52 932 92 934
rect 52 924 92 926
rect 208 911 248 913
rect 1716 911 1756 913
rect 208 903 248 905
rect 1716 903 1756 905
rect 1882 874 1922 876
rect 1882 866 1922 868
rect 1560 846 1600 848
rect 1560 838 1600 840
rect 180 822 220 824
rect 180 814 220 816
rect 517 813 519 833
rect 1716 825 1756 827
rect 1716 817 1756 819
rect 215 646 255 648
rect 215 638 255 640
rect 1716 636 1756 638
rect 1716 628 1756 630
rect 381 609 421 611
rect 381 601 421 603
rect 1882 599 1922 601
rect 1882 591 1922 593
rect 59 581 99 583
rect 923 576 963 578
rect 59 573 99 575
rect 1560 571 1600 573
rect 923 568 963 570
rect 1560 563 1600 565
rect 215 560 255 562
rect 215 552 255 554
rect 1716 550 1756 552
rect 1716 542 1756 544
rect 1147 511 1187 513
rect 1147 503 1187 505
rect 187 471 227 473
rect 187 463 227 465
rect 520 462 522 482
rect 1718 442 1758 444
rect 1718 434 1758 436
rect 1884 405 1924 407
rect 1884 397 1924 399
rect 1562 377 1602 379
rect 920 369 980 371
rect 1562 369 1602 371
rect 920 361 980 363
rect 1718 356 1758 358
rect 920 353 980 355
rect 1718 348 1758 350
rect 1109 328 1169 330
rect 1109 320 1169 322
rect 1109 312 1169 314
rect 185 305 225 307
rect 185 297 225 299
rect 926 285 966 287
rect 926 277 966 279
rect 351 268 391 270
rect 351 260 391 262
rect 29 240 69 242
rect 1725 241 1765 243
rect 29 232 69 234
rect 1725 233 1765 235
rect 185 219 225 221
rect 185 211 225 213
rect 912 203 992 205
rect 1891 204 1931 206
rect 912 195 992 197
rect 1891 196 1931 198
rect 912 187 992 189
rect 912 179 992 181
rect 1569 176 1609 178
rect 1569 168 1609 170
rect 1131 154 1211 156
rect 1725 155 1765 157
rect 1131 146 1211 148
rect 1725 147 1765 149
rect 157 130 197 132
rect 157 122 197 124
rect 499 121 501 141
rect 1131 138 1211 140
rect 1131 130 1211 132
rect 916 106 976 108
rect 916 98 976 100
rect 916 90 976 92
rect 922 33 962 35
rect 922 25 962 27
rect 184 -37 224 -35
rect 184 -45 224 -43
rect 350 -74 390 -72
rect 350 -82 390 -80
rect 28 -102 68 -100
rect 28 -110 68 -108
rect 184 -123 224 -121
rect 184 -131 224 -129
rect 156 -212 196 -210
rect 156 -220 196 -218
rect 493 -221 495 -201
rect 880 -303 960 -301
rect 880 -311 960 -309
rect 178 -319 218 -317
rect 880 -319 960 -317
rect 178 -327 218 -325
rect 880 -327 960 -325
rect 880 -335 960 -333
rect 344 -356 384 -354
rect 344 -364 384 -362
rect 22 -384 62 -382
rect 1164 -388 1244 -386
rect 22 -392 62 -390
rect 1164 -396 1244 -394
rect 178 -405 218 -403
rect 1164 -404 1244 -402
rect 178 -413 218 -411
rect 1164 -412 1244 -410
rect 1164 -420 1244 -418
rect 902 -464 982 -462
rect 902 -472 982 -470
rect 902 -480 982 -478
rect 902 -488 982 -486
rect 150 -494 190 -492
rect 150 -502 190 -500
rect 909 -608 969 -606
rect 909 -616 969 -614
rect 909 -624 969 -622
rect 926 -698 966 -696
rect 926 -706 966 -704
<< ptransistor >>
rect 153 997 193 999
rect 153 989 193 991
rect 319 960 359 962
rect 319 952 359 954
rect -3 932 37 934
rect -3 924 37 926
rect 153 911 193 913
rect 1661 911 1701 913
rect 153 903 193 905
rect 1661 903 1701 905
rect 517 847 519 887
rect 1827 874 1867 876
rect 1827 866 1867 868
rect 1505 846 1545 848
rect 1505 838 1545 840
rect 125 822 165 824
rect 125 814 165 816
rect 1661 825 1701 827
rect 1661 817 1701 819
rect 160 646 200 648
rect 160 638 200 640
rect 1661 636 1701 638
rect 1661 628 1701 630
rect 326 609 366 611
rect 326 601 366 603
rect 1827 599 1867 601
rect 1827 591 1867 593
rect 4 581 44 583
rect 868 576 908 578
rect 4 573 44 575
rect 1505 571 1545 573
rect 868 568 908 570
rect 1505 563 1545 565
rect 160 560 200 562
rect 160 552 200 554
rect 1661 550 1701 552
rect 1661 542 1701 544
rect 520 496 522 536
rect 1092 511 1132 513
rect 1092 503 1132 505
rect 132 471 172 473
rect 132 463 172 465
rect 1663 442 1703 444
rect 1663 434 1703 436
rect 1829 405 1869 407
rect 1829 397 1869 399
rect 1507 377 1547 379
rect 862 369 902 371
rect 1507 369 1547 371
rect 862 361 902 363
rect 1663 356 1703 358
rect 862 353 902 355
rect 1663 348 1703 350
rect 1051 328 1091 330
rect 1051 320 1091 322
rect 1051 312 1091 314
rect 130 305 170 307
rect 130 297 170 299
rect 871 285 911 287
rect 871 277 911 279
rect 296 268 336 270
rect 296 260 336 262
rect -26 240 14 242
rect 1670 241 1710 243
rect -26 232 14 234
rect 1670 233 1710 235
rect 130 219 170 221
rect 130 211 170 213
rect 848 203 888 205
rect 1836 204 1876 206
rect 499 155 501 195
rect 848 195 888 197
rect 1836 196 1876 198
rect 848 187 888 189
rect 848 179 888 181
rect 1514 176 1554 178
rect 1514 168 1554 170
rect 1067 154 1107 156
rect 1670 155 1710 157
rect 1067 146 1107 148
rect 1670 147 1710 149
rect 102 130 142 132
rect 102 122 142 124
rect 1067 138 1107 140
rect 1067 130 1107 132
rect 858 106 898 108
rect 858 98 898 100
rect 858 90 898 92
rect 867 33 907 35
rect 867 25 907 27
rect 129 -37 169 -35
rect 129 -45 169 -43
rect 295 -74 335 -72
rect 295 -82 335 -80
rect -27 -102 13 -100
rect -27 -110 13 -108
rect 129 -123 169 -121
rect 129 -131 169 -129
rect 493 -187 495 -147
rect 101 -212 141 -210
rect 101 -220 141 -218
rect 816 -303 856 -301
rect 816 -311 856 -309
rect 123 -319 163 -317
rect 816 -319 856 -317
rect 123 -327 163 -325
rect 816 -327 856 -325
rect 816 -335 856 -333
rect 289 -356 329 -354
rect 289 -364 329 -362
rect -33 -384 7 -382
rect 1100 -388 1140 -386
rect -33 -392 7 -390
rect 1100 -396 1140 -394
rect 123 -405 163 -403
rect 1100 -404 1140 -402
rect 123 -413 163 -411
rect 1100 -412 1140 -410
rect 1100 -420 1140 -418
rect 838 -464 878 -462
rect 838 -472 878 -470
rect 838 -480 878 -478
rect 838 -488 878 -486
rect 95 -494 135 -492
rect 95 -502 135 -500
rect 851 -608 891 -606
rect 851 -616 891 -614
rect 851 -624 891 -622
rect 871 -698 911 -696
rect 871 -706 911 -704
<< ndiffusion >>
rect 208 999 248 1000
rect 208 996 248 997
rect 208 991 248 992
rect 208 988 248 989
rect 374 962 414 963
rect 374 959 414 960
rect 374 954 414 955
rect 374 951 414 952
rect 52 934 92 935
rect 52 931 92 932
rect 52 926 92 927
rect 52 923 92 924
rect 208 913 248 914
rect 208 910 248 911
rect 1716 913 1756 914
rect 208 905 248 906
rect 208 902 248 903
rect 1716 910 1756 911
rect 1716 905 1756 906
rect 1716 902 1756 903
rect 1882 876 1922 877
rect 1882 873 1922 874
rect 1882 868 1922 869
rect 1882 865 1922 866
rect 1560 848 1600 849
rect 1560 845 1600 846
rect 1560 840 1600 841
rect 1560 837 1600 838
rect 180 824 220 825
rect 180 821 220 822
rect 180 816 220 817
rect 180 813 220 814
rect 516 813 517 833
rect 519 813 520 833
rect 1716 827 1756 828
rect 1716 824 1756 825
rect 1716 819 1756 820
rect 1716 816 1756 817
rect 215 648 255 649
rect 215 645 255 646
rect 215 640 255 641
rect 215 637 255 638
rect 1716 638 1756 639
rect 1716 635 1756 636
rect 1716 630 1756 631
rect 1716 627 1756 628
rect 381 611 421 612
rect 381 608 421 609
rect 381 603 421 604
rect 381 600 421 601
rect 1882 601 1922 602
rect 1882 598 1922 599
rect 1882 593 1922 594
rect 1882 590 1922 591
rect 59 583 99 584
rect 59 580 99 581
rect 59 575 99 576
rect 923 578 963 579
rect 59 572 99 573
rect 923 575 963 576
rect 923 570 963 571
rect 1560 573 1600 574
rect 923 567 963 568
rect 215 562 255 563
rect 1560 570 1600 571
rect 1560 565 1600 566
rect 215 559 255 560
rect 1560 562 1600 563
rect 215 554 255 555
rect 215 551 255 552
rect 1716 552 1756 553
rect 1716 549 1756 550
rect 1716 544 1756 545
rect 1716 541 1756 542
rect 1147 513 1187 514
rect 1147 510 1187 511
rect 1147 505 1187 506
rect 1147 502 1187 503
rect 187 473 227 474
rect 187 470 227 471
rect 187 465 227 466
rect 187 462 227 463
rect 519 462 520 482
rect 522 462 523 482
rect 1718 444 1758 445
rect 1718 441 1758 442
rect 1718 436 1758 437
rect 1718 433 1758 434
rect 1884 407 1924 408
rect 1884 404 1924 405
rect 1884 399 1924 400
rect 1884 396 1924 397
rect 1562 379 1602 380
rect 920 371 980 372
rect 920 368 980 369
rect 1562 376 1602 377
rect 1562 371 1602 372
rect 1562 368 1602 369
rect 920 363 980 364
rect 920 360 980 361
rect 920 355 980 356
rect 1718 358 1758 359
rect 920 352 980 353
rect 1718 355 1758 356
rect 1718 350 1758 351
rect 1718 347 1758 348
rect 1109 330 1169 331
rect 1109 327 1169 328
rect 1109 322 1169 323
rect 1109 319 1169 320
rect 1109 314 1169 315
rect 185 307 225 308
rect 1109 311 1169 312
rect 185 304 225 305
rect 185 299 225 300
rect 185 296 225 297
rect 926 287 966 288
rect 926 284 966 285
rect 926 279 966 280
rect 926 276 966 277
rect 351 270 391 271
rect 351 267 391 268
rect 351 262 391 263
rect 351 259 391 260
rect 29 242 69 243
rect 1725 243 1765 244
rect 29 239 69 240
rect 29 234 69 235
rect 1725 240 1765 241
rect 1725 235 1765 236
rect 29 231 69 232
rect 1725 232 1765 233
rect 185 221 225 222
rect 185 218 225 219
rect 185 213 225 214
rect 185 210 225 211
rect 912 205 992 206
rect 1891 206 1931 207
rect 912 202 992 203
rect 912 197 992 198
rect 1891 203 1931 204
rect 1891 198 1931 199
rect 912 194 992 195
rect 1891 195 1931 196
rect 912 189 992 190
rect 912 186 992 187
rect 912 181 992 182
rect 912 178 992 179
rect 1569 178 1609 179
rect 1569 175 1609 176
rect 1569 170 1609 171
rect 1569 167 1609 168
rect 1131 156 1211 157
rect 1725 157 1765 158
rect 1131 153 1211 154
rect 1131 148 1211 149
rect 1725 154 1765 155
rect 1725 149 1765 150
rect 157 132 197 133
rect 157 129 197 130
rect 157 124 197 125
rect 157 121 197 122
rect 498 121 499 141
rect 501 121 502 141
rect 1131 145 1211 146
rect 1725 146 1765 147
rect 1131 140 1211 141
rect 1131 137 1211 138
rect 1131 132 1211 133
rect 1131 129 1211 130
rect 916 108 976 109
rect 916 105 976 106
rect 916 100 976 101
rect 916 97 976 98
rect 916 92 976 93
rect 916 89 976 90
rect 922 35 962 36
rect 922 32 962 33
rect 922 27 962 28
rect 922 24 962 25
rect 184 -35 224 -34
rect 184 -38 224 -37
rect 184 -43 224 -42
rect 184 -46 224 -45
rect 350 -72 390 -71
rect 350 -75 390 -74
rect 350 -80 390 -79
rect 350 -83 390 -82
rect 28 -100 68 -99
rect 28 -103 68 -102
rect 28 -108 68 -107
rect 28 -111 68 -110
rect 184 -121 224 -120
rect 184 -124 224 -123
rect 184 -129 224 -128
rect 184 -132 224 -131
rect 156 -210 196 -209
rect 156 -213 196 -212
rect 156 -218 196 -217
rect 156 -221 196 -220
rect 492 -221 493 -201
rect 495 -221 496 -201
rect 880 -301 960 -300
rect 880 -304 960 -303
rect 880 -309 960 -308
rect 178 -317 218 -316
rect 178 -320 218 -319
rect 880 -312 960 -311
rect 880 -317 960 -316
rect 178 -325 218 -324
rect 178 -328 218 -327
rect 880 -320 960 -319
rect 880 -325 960 -324
rect 880 -328 960 -327
rect 880 -333 960 -332
rect 880 -336 960 -335
rect 344 -354 384 -353
rect 344 -357 384 -356
rect 344 -362 384 -361
rect 344 -365 384 -364
rect 22 -382 62 -381
rect 22 -385 62 -384
rect 1164 -386 1244 -385
rect 22 -390 62 -389
rect 22 -393 62 -392
rect 1164 -389 1244 -388
rect 1164 -394 1244 -393
rect 178 -403 218 -402
rect 1164 -397 1244 -396
rect 1164 -402 1244 -401
rect 178 -406 218 -405
rect 178 -411 218 -410
rect 1164 -405 1244 -404
rect 1164 -410 1244 -409
rect 178 -414 218 -413
rect 1164 -413 1244 -412
rect 1164 -418 1244 -417
rect 1164 -421 1244 -420
rect 902 -462 982 -461
rect 902 -465 982 -464
rect 902 -470 982 -469
rect 902 -473 982 -472
rect 902 -478 982 -477
rect 902 -481 982 -480
rect 902 -486 982 -485
rect 150 -492 190 -491
rect 902 -489 982 -488
rect 150 -495 190 -494
rect 150 -500 190 -499
rect 150 -503 190 -502
rect 909 -606 969 -605
rect 909 -609 969 -608
rect 909 -614 969 -613
rect 909 -617 969 -616
rect 909 -622 969 -621
rect 909 -625 969 -624
rect 926 -696 966 -695
rect 926 -699 966 -698
rect 926 -704 966 -703
rect 926 -707 966 -706
<< pdiffusion >>
rect 153 999 193 1000
rect 153 996 193 997
rect 153 991 193 992
rect 153 988 193 989
rect 319 962 359 963
rect 319 959 359 960
rect 319 954 359 955
rect 319 951 359 952
rect -3 934 37 935
rect -3 931 37 932
rect -3 926 37 927
rect -3 923 37 924
rect 153 913 193 914
rect 153 910 193 911
rect 153 905 193 906
rect 1661 913 1701 914
rect 1661 910 1701 911
rect 153 902 193 903
rect 1661 905 1701 906
rect 1661 902 1701 903
rect 516 847 517 887
rect 519 847 520 887
rect 1827 876 1867 877
rect 1827 873 1867 874
rect 1827 868 1867 869
rect 1827 865 1867 866
rect 1505 848 1545 849
rect 1505 845 1545 846
rect 1505 840 1545 841
rect 1505 837 1545 838
rect 125 824 165 825
rect 125 821 165 822
rect 125 816 165 817
rect 125 813 165 814
rect 1661 827 1701 828
rect 1661 824 1701 825
rect 1661 819 1701 820
rect 1661 816 1701 817
rect 160 648 200 649
rect 160 645 200 646
rect 160 640 200 641
rect 160 637 200 638
rect 1661 638 1701 639
rect 1661 635 1701 636
rect 1661 630 1701 631
rect 1661 627 1701 628
rect 326 611 366 612
rect 326 608 366 609
rect 326 603 366 604
rect 326 600 366 601
rect 1827 601 1867 602
rect 1827 598 1867 599
rect 1827 593 1867 594
rect 1827 590 1867 591
rect 4 583 44 584
rect 4 580 44 581
rect 4 575 44 576
rect 868 578 908 579
rect 868 575 908 576
rect 4 572 44 573
rect 868 570 908 571
rect 1505 573 1545 574
rect 1505 570 1545 571
rect 868 567 908 568
rect 160 562 200 563
rect 1505 565 1545 566
rect 1505 562 1545 563
rect 160 559 200 560
rect 160 554 200 555
rect 160 551 200 552
rect 1661 552 1701 553
rect 1661 549 1701 550
rect 1661 544 1701 545
rect 1661 541 1701 542
rect 519 496 520 536
rect 522 496 523 536
rect 1092 513 1132 514
rect 1092 510 1132 511
rect 1092 505 1132 506
rect 1092 502 1132 503
rect 132 473 172 474
rect 132 470 172 471
rect 132 465 172 466
rect 132 462 172 463
rect 1663 444 1703 445
rect 1663 441 1703 442
rect 1663 436 1703 437
rect 1663 433 1703 434
rect 1829 407 1869 408
rect 1829 404 1869 405
rect 1829 399 1869 400
rect 1829 396 1869 397
rect 1507 379 1547 380
rect 1507 376 1547 377
rect 862 371 902 372
rect 862 368 902 369
rect 862 363 902 364
rect 1507 371 1547 372
rect 1507 368 1547 369
rect 862 360 902 361
rect 862 355 902 356
rect 1663 358 1703 359
rect 1663 355 1703 356
rect 862 352 902 353
rect 1663 350 1703 351
rect 1663 347 1703 348
rect 1051 330 1091 331
rect 1051 327 1091 328
rect 1051 322 1091 323
rect 1051 319 1091 320
rect 130 307 170 308
rect 1051 314 1091 315
rect 1051 311 1091 312
rect 130 304 170 305
rect 130 299 170 300
rect 130 296 170 297
rect 871 287 911 288
rect 871 284 911 285
rect 871 279 911 280
rect 871 276 911 277
rect 296 270 336 271
rect 296 267 336 268
rect 296 262 336 263
rect 296 259 336 260
rect -26 242 14 243
rect 1670 243 1710 244
rect 1670 240 1710 241
rect -26 239 14 240
rect -26 234 14 235
rect 1670 235 1710 236
rect 1670 232 1710 233
rect -26 231 14 232
rect 130 221 170 222
rect 130 218 170 219
rect 130 213 170 214
rect 130 210 170 211
rect 848 205 888 206
rect 1836 206 1876 207
rect 1836 203 1876 204
rect 848 202 888 203
rect 498 155 499 195
rect 501 155 502 195
rect 848 197 888 198
rect 1836 198 1876 199
rect 1836 195 1876 196
rect 848 194 888 195
rect 848 189 888 190
rect 848 186 888 187
rect 848 181 888 182
rect 848 178 888 179
rect 1514 178 1554 179
rect 1514 175 1554 176
rect 1514 170 1554 171
rect 1514 167 1554 168
rect 1067 156 1107 157
rect 1670 157 1710 158
rect 1670 154 1710 155
rect 1067 153 1107 154
rect 1067 148 1107 149
rect 1670 149 1710 150
rect 1670 146 1710 147
rect 1067 145 1107 146
rect 102 132 142 133
rect 102 129 142 130
rect 102 124 142 125
rect 102 121 142 122
rect 1067 140 1107 141
rect 1067 137 1107 138
rect 1067 132 1107 133
rect 1067 129 1107 130
rect 858 108 898 109
rect 858 105 898 106
rect 858 100 898 101
rect 858 97 898 98
rect 858 92 898 93
rect 858 89 898 90
rect 867 35 907 36
rect 867 32 907 33
rect 867 27 907 28
rect 867 24 907 25
rect 129 -35 169 -34
rect 129 -38 169 -37
rect 129 -43 169 -42
rect 129 -46 169 -45
rect 295 -72 335 -71
rect 295 -75 335 -74
rect 295 -80 335 -79
rect 295 -83 335 -82
rect -27 -100 13 -99
rect -27 -103 13 -102
rect -27 -108 13 -107
rect -27 -111 13 -110
rect 129 -121 169 -120
rect 129 -124 169 -123
rect 129 -129 169 -128
rect 129 -132 169 -131
rect 492 -187 493 -147
rect 495 -187 496 -147
rect 101 -210 141 -209
rect 101 -213 141 -212
rect 101 -218 141 -217
rect 101 -221 141 -220
rect 816 -301 856 -300
rect 816 -304 856 -303
rect 816 -309 856 -308
rect 816 -312 856 -311
rect 123 -317 163 -316
rect 123 -320 163 -319
rect 123 -325 163 -324
rect 816 -317 856 -316
rect 816 -320 856 -319
rect 123 -328 163 -327
rect 816 -325 856 -324
rect 816 -328 856 -327
rect 816 -333 856 -332
rect 816 -336 856 -335
rect 289 -354 329 -353
rect 289 -357 329 -356
rect 289 -362 329 -361
rect 289 -365 329 -364
rect -33 -382 7 -381
rect -33 -385 7 -384
rect -33 -390 7 -389
rect 1100 -386 1140 -385
rect 1100 -389 1140 -388
rect -33 -393 7 -392
rect 1100 -394 1140 -393
rect 1100 -397 1140 -396
rect 123 -403 163 -402
rect 1100 -402 1140 -401
rect 1100 -405 1140 -404
rect 123 -406 163 -405
rect 123 -411 163 -410
rect 1100 -410 1140 -409
rect 1100 -413 1140 -412
rect 123 -414 163 -413
rect 1100 -418 1140 -417
rect 1100 -421 1140 -420
rect 838 -462 878 -461
rect 838 -465 878 -464
rect 838 -470 878 -469
rect 838 -473 878 -472
rect 838 -478 878 -477
rect 838 -481 878 -480
rect 95 -492 135 -491
rect 838 -486 878 -485
rect 838 -489 878 -488
rect 95 -495 135 -494
rect 95 -500 135 -499
rect 95 -503 135 -502
rect 851 -606 891 -605
rect 851 -609 891 -608
rect 851 -614 891 -613
rect 851 -617 891 -616
rect 851 -622 891 -621
rect 851 -625 891 -624
rect 871 -696 911 -695
rect 871 -699 911 -698
rect 871 -704 911 -703
rect 871 -707 911 -706
<< ndcontact >>
rect 208 1000 248 1004
rect 208 992 248 996
rect 208 984 248 988
rect 374 963 414 967
rect 374 955 414 959
rect 374 947 414 951
rect 52 935 92 939
rect 52 927 92 931
rect 52 919 92 923
rect 208 914 248 918
rect 1716 914 1756 918
rect 208 906 248 910
rect 1716 906 1756 910
rect 208 898 248 902
rect 1716 898 1756 902
rect 1882 877 1922 881
rect 1882 869 1922 873
rect 1882 861 1922 865
rect 1560 849 1600 853
rect 1560 841 1600 845
rect 1560 833 1600 837
rect 180 825 220 829
rect 180 817 220 821
rect 512 813 516 833
rect 520 813 524 833
rect 1716 828 1756 832
rect 1716 820 1756 824
rect 180 809 220 813
rect 1716 812 1756 816
rect 215 649 255 653
rect 215 641 255 645
rect 215 633 255 637
rect 1716 639 1756 643
rect 1716 631 1756 635
rect 1716 623 1756 627
rect 381 612 421 616
rect 381 604 421 608
rect 381 596 421 600
rect 1882 602 1922 606
rect 1882 594 1922 598
rect 59 584 99 588
rect 1882 586 1922 590
rect 59 576 99 580
rect 923 579 963 583
rect 59 568 99 572
rect 923 571 963 575
rect 1560 574 1600 578
rect 215 563 255 567
rect 923 563 963 567
rect 1560 566 1600 570
rect 215 555 255 559
rect 1560 558 1600 562
rect 215 547 255 551
rect 1716 553 1756 557
rect 1716 545 1756 549
rect 1716 537 1756 541
rect 1147 514 1187 518
rect 1147 506 1187 510
rect 1147 498 1187 502
rect 187 474 227 478
rect 187 466 227 470
rect 515 462 519 482
rect 523 462 527 482
rect 187 458 227 462
rect 1718 445 1758 449
rect 1718 437 1758 441
rect 1718 429 1758 433
rect 1884 408 1924 412
rect 1884 400 1924 404
rect 1884 392 1924 396
rect 1562 380 1602 384
rect 920 372 980 376
rect 1562 372 1602 376
rect 920 364 980 368
rect 1562 364 1602 368
rect 920 356 980 360
rect 1718 359 1758 363
rect 920 348 980 352
rect 1718 351 1758 355
rect 1718 343 1758 347
rect 1109 331 1169 335
rect 1109 323 1169 327
rect 185 308 225 312
rect 1109 315 1169 319
rect 1109 307 1169 311
rect 185 300 225 304
rect 185 292 225 296
rect 926 288 966 292
rect 926 280 966 284
rect 351 271 391 275
rect 926 272 966 276
rect 351 263 391 267
rect 351 255 391 259
rect 29 243 69 247
rect 1725 244 1765 248
rect 29 235 69 239
rect 1725 236 1765 240
rect 29 227 69 231
rect 1725 228 1765 232
rect 185 222 225 226
rect 185 214 225 218
rect 185 206 225 210
rect 912 206 992 210
rect 1891 207 1931 211
rect 912 198 992 202
rect 1891 199 1931 203
rect 912 190 992 194
rect 1891 191 1931 195
rect 912 182 992 186
rect 912 174 992 178
rect 1569 179 1609 183
rect 1569 171 1609 175
rect 1569 163 1609 167
rect 1131 157 1211 161
rect 1725 158 1765 162
rect 1131 149 1211 153
rect 1725 150 1765 154
rect 157 133 197 137
rect 157 125 197 129
rect 494 121 498 141
rect 502 121 506 141
rect 1131 141 1211 145
rect 1725 142 1765 146
rect 1131 133 1211 137
rect 1131 125 1211 129
rect 157 117 197 121
rect 916 109 976 113
rect 916 101 976 105
rect 916 93 976 97
rect 916 85 976 89
rect 922 36 962 40
rect 922 28 962 32
rect 922 20 962 24
rect 184 -34 224 -30
rect 184 -42 224 -38
rect 184 -50 224 -46
rect 350 -71 390 -67
rect 350 -79 390 -75
rect 350 -87 390 -83
rect 28 -99 68 -95
rect 28 -107 68 -103
rect 28 -115 68 -111
rect 184 -120 224 -116
rect 184 -128 224 -124
rect 184 -136 224 -132
rect 156 -209 196 -205
rect 156 -217 196 -213
rect 488 -221 492 -201
rect 496 -221 500 -201
rect 156 -225 196 -221
rect 880 -300 960 -296
rect 880 -308 960 -304
rect 178 -316 218 -312
rect 880 -316 960 -312
rect 178 -324 218 -320
rect 880 -324 960 -320
rect 178 -332 218 -328
rect 880 -332 960 -328
rect 880 -340 960 -336
rect 344 -353 384 -349
rect 344 -361 384 -357
rect 344 -369 384 -365
rect 22 -381 62 -377
rect 22 -389 62 -385
rect 1164 -385 1244 -381
rect 22 -397 62 -393
rect 1164 -393 1244 -389
rect 178 -402 218 -398
rect 1164 -401 1244 -397
rect 178 -410 218 -406
rect 1164 -409 1244 -405
rect 178 -418 218 -414
rect 1164 -417 1244 -413
rect 1164 -425 1244 -421
rect 902 -461 982 -457
rect 902 -469 982 -465
rect 902 -477 982 -473
rect 150 -491 190 -487
rect 902 -485 982 -481
rect 902 -493 982 -489
rect 150 -499 190 -495
rect 150 -507 190 -503
rect 909 -605 969 -601
rect 909 -613 969 -609
rect 909 -621 969 -617
rect 909 -629 969 -625
rect 926 -695 966 -691
rect 926 -703 966 -699
rect 926 -711 966 -707
<< pdcontact >>
rect 153 1000 193 1004
rect 153 992 193 996
rect 153 984 193 988
rect 319 963 359 967
rect 319 955 359 959
rect 319 947 359 951
rect -3 935 37 939
rect -3 927 37 931
rect -3 919 37 923
rect 153 914 193 918
rect 1661 914 1701 918
rect 153 906 193 910
rect 1661 906 1701 910
rect 153 898 193 902
rect 1661 898 1701 902
rect 512 847 516 887
rect 520 847 524 887
rect 1827 877 1867 881
rect 1827 869 1867 873
rect 1827 861 1867 865
rect 1505 849 1545 853
rect 1505 841 1545 845
rect 1505 833 1545 837
rect 125 825 165 829
rect 125 817 165 821
rect 125 809 165 813
rect 1661 828 1701 832
rect 1661 820 1701 824
rect 1661 812 1701 816
rect 160 649 200 653
rect 160 641 200 645
rect 1661 639 1701 643
rect 160 633 200 637
rect 1661 631 1701 635
rect 1661 623 1701 627
rect 326 612 366 616
rect 326 604 366 608
rect 1827 602 1867 606
rect 326 596 366 600
rect 1827 594 1867 598
rect 4 584 44 588
rect 1827 586 1867 590
rect 4 576 44 580
rect 868 579 908 583
rect 4 568 44 572
rect 868 571 908 575
rect 1505 574 1545 578
rect 160 563 200 567
rect 868 563 908 567
rect 1505 566 1545 570
rect 160 555 200 559
rect 1505 558 1545 562
rect 1661 553 1701 557
rect 160 547 200 551
rect 1661 545 1701 549
rect 1661 537 1701 541
rect 515 496 519 536
rect 523 496 527 536
rect 1092 514 1132 518
rect 1092 506 1132 510
rect 1092 498 1132 502
rect 132 474 172 478
rect 132 466 172 470
rect 132 458 172 462
rect 1663 445 1703 449
rect 1663 437 1703 441
rect 1663 429 1703 433
rect 1829 408 1869 412
rect 1829 400 1869 404
rect 1829 392 1869 396
rect 1507 380 1547 384
rect 862 372 902 376
rect 1507 372 1547 376
rect 862 364 902 368
rect 1507 364 1547 368
rect 862 356 902 360
rect 1663 359 1703 363
rect 862 348 902 352
rect 1663 351 1703 355
rect 1663 343 1703 347
rect 1051 331 1091 335
rect 1051 323 1091 327
rect 1051 315 1091 319
rect 130 308 170 312
rect 1051 307 1091 311
rect 130 300 170 304
rect 130 292 170 296
rect 871 288 911 292
rect 871 280 911 284
rect 296 271 336 275
rect 871 272 911 276
rect 296 263 336 267
rect 296 255 336 259
rect -26 243 14 247
rect 1670 244 1710 248
rect -26 235 14 239
rect 1670 236 1710 240
rect -26 227 14 231
rect 1670 228 1710 232
rect 130 222 170 226
rect 130 214 170 218
rect 130 206 170 210
rect 848 206 888 210
rect 1836 207 1876 211
rect 848 198 888 202
rect 494 155 498 195
rect 502 155 506 195
rect 1836 199 1876 203
rect 848 190 888 194
rect 1836 191 1876 195
rect 848 182 888 186
rect 1514 179 1554 183
rect 848 174 888 178
rect 1514 171 1554 175
rect 1514 163 1554 167
rect 1067 157 1107 161
rect 1670 158 1710 162
rect 1067 149 1107 153
rect 1670 150 1710 154
rect 1067 141 1107 145
rect 102 133 142 137
rect 102 125 142 129
rect 102 117 142 121
rect 1670 142 1710 146
rect 1067 133 1107 137
rect 1067 125 1107 129
rect 858 109 898 113
rect 858 101 898 105
rect 858 93 898 97
rect 858 85 898 89
rect 867 36 907 40
rect 867 28 907 32
rect 867 20 907 24
rect 129 -34 169 -30
rect 129 -42 169 -38
rect 129 -50 169 -46
rect 295 -71 335 -67
rect 295 -79 335 -75
rect 295 -87 335 -83
rect -27 -99 13 -95
rect -27 -107 13 -103
rect -27 -115 13 -111
rect 129 -120 169 -116
rect 129 -128 169 -124
rect 129 -136 169 -132
rect 488 -187 492 -147
rect 496 -187 500 -147
rect 101 -209 141 -205
rect 101 -217 141 -213
rect 101 -225 141 -221
rect 816 -300 856 -296
rect 816 -308 856 -304
rect 123 -316 163 -312
rect 816 -316 856 -312
rect 123 -324 163 -320
rect 816 -324 856 -320
rect 123 -332 163 -328
rect 816 -332 856 -328
rect 816 -340 856 -336
rect 289 -353 329 -349
rect 289 -361 329 -357
rect 289 -369 329 -365
rect -33 -381 7 -377
rect -33 -389 7 -385
rect 1100 -385 1140 -381
rect -33 -397 7 -393
rect 1100 -393 1140 -389
rect 123 -402 163 -398
rect 1100 -401 1140 -397
rect 123 -410 163 -406
rect 1100 -409 1140 -405
rect 123 -418 163 -414
rect 1100 -417 1140 -413
rect 1100 -425 1140 -421
rect 838 -461 878 -457
rect 838 -469 878 -465
rect 838 -477 878 -473
rect 838 -485 878 -481
rect 95 -491 135 -487
rect 838 -493 878 -489
rect 95 -499 135 -495
rect 95 -507 135 -503
rect 851 -605 891 -601
rect 851 -613 891 -609
rect 851 -621 891 -617
rect 851 -629 891 -625
rect 871 -695 911 -691
rect 871 -703 911 -699
rect 871 -711 911 -707
<< polysilicon >>
rect 142 997 153 999
rect 193 997 208 999
rect 248 997 252 999
rect 142 989 153 991
rect 193 989 208 991
rect 248 989 252 991
rect 308 960 319 962
rect 359 960 374 962
rect 414 960 418 962
rect 308 952 319 954
rect 359 952 374 954
rect 414 952 418 954
rect -14 932 -3 934
rect 37 932 52 934
rect 92 932 96 934
rect -14 924 -3 926
rect 37 924 52 926
rect 92 924 96 926
rect 142 911 153 913
rect 193 911 208 913
rect 248 911 252 913
rect 1650 911 1661 913
rect 1701 911 1716 913
rect 1756 911 1760 913
rect 142 903 153 905
rect 193 903 208 905
rect 248 903 252 905
rect 1650 903 1661 905
rect 1701 903 1716 905
rect 1756 903 1760 905
rect 517 887 519 890
rect 1816 874 1827 876
rect 1867 874 1882 876
rect 1922 874 1926 876
rect 1816 866 1827 868
rect 1867 866 1882 868
rect 1922 866 1926 868
rect 517 833 519 847
rect 1494 846 1505 848
rect 1545 846 1560 848
rect 1600 846 1604 848
rect 1494 838 1505 840
rect 1545 838 1560 840
rect 1600 838 1604 840
rect 114 822 125 824
rect 165 822 180 824
rect 220 822 224 824
rect 114 814 125 816
rect 165 814 180 816
rect 220 814 224 816
rect 1650 825 1661 827
rect 1701 825 1716 827
rect 1756 825 1760 827
rect 1650 817 1661 819
rect 1701 817 1716 819
rect 1756 817 1760 819
rect 517 810 519 813
rect 149 646 160 648
rect 200 646 215 648
rect 255 646 259 648
rect 149 638 160 640
rect 200 638 215 640
rect 255 638 259 640
rect 1650 636 1661 638
rect 1701 636 1716 638
rect 1756 636 1760 638
rect 1650 628 1661 630
rect 1701 628 1716 630
rect 1756 628 1760 630
rect 315 609 326 611
rect 366 609 381 611
rect 421 609 425 611
rect 315 601 326 603
rect 366 601 381 603
rect 421 601 425 603
rect 1816 599 1827 601
rect 1867 599 1882 601
rect 1922 599 1926 601
rect 1816 591 1827 593
rect 1867 591 1882 593
rect 1922 591 1926 593
rect -7 581 4 583
rect 44 581 59 583
rect 99 581 103 583
rect 857 576 868 578
rect 908 576 923 578
rect 963 576 967 578
rect -7 573 4 575
rect 44 573 59 575
rect 99 573 103 575
rect 1494 571 1505 573
rect 1545 571 1560 573
rect 1600 571 1604 573
rect 857 568 868 570
rect 908 568 923 570
rect 963 568 967 570
rect 1494 563 1505 565
rect 1545 563 1560 565
rect 1600 563 1604 565
rect 149 560 160 562
rect 200 560 215 562
rect 255 560 259 562
rect 149 552 160 554
rect 200 552 215 554
rect 255 552 259 554
rect 1650 550 1661 552
rect 1701 550 1716 552
rect 1756 550 1760 552
rect 1650 542 1661 544
rect 1701 542 1716 544
rect 1756 542 1760 544
rect 520 536 522 539
rect 1081 511 1092 513
rect 1132 511 1147 513
rect 1187 511 1191 513
rect 1081 503 1092 505
rect 1132 503 1147 505
rect 1187 503 1191 505
rect 520 482 522 496
rect 121 471 132 473
rect 172 471 187 473
rect 227 471 231 473
rect 121 463 132 465
rect 172 463 187 465
rect 227 463 231 465
rect 520 459 522 462
rect 1652 442 1663 444
rect 1703 442 1718 444
rect 1758 442 1762 444
rect 1652 434 1663 436
rect 1703 434 1718 436
rect 1758 434 1762 436
rect 1818 405 1829 407
rect 1869 405 1884 407
rect 1924 405 1928 407
rect 1818 397 1829 399
rect 1869 397 1884 399
rect 1924 397 1928 399
rect 1496 377 1507 379
rect 1547 377 1562 379
rect 1602 377 1606 379
rect 851 369 862 371
rect 902 369 920 371
rect 980 369 985 371
rect 1496 369 1507 371
rect 1547 369 1562 371
rect 1602 369 1606 371
rect 851 361 862 363
rect 902 361 920 363
rect 980 361 985 363
rect 1652 356 1663 358
rect 1703 356 1718 358
rect 1758 356 1762 358
rect 851 353 862 355
rect 902 353 920 355
rect 980 353 985 355
rect 1652 348 1663 350
rect 1703 348 1718 350
rect 1758 348 1762 350
rect 1040 328 1051 330
rect 1091 328 1109 330
rect 1169 328 1174 330
rect 1040 320 1051 322
rect 1091 320 1109 322
rect 1169 320 1174 322
rect 1040 312 1051 314
rect 1091 312 1109 314
rect 1169 312 1174 314
rect 119 305 130 307
rect 170 305 185 307
rect 225 305 229 307
rect 119 297 130 299
rect 170 297 185 299
rect 225 297 229 299
rect 860 285 871 287
rect 911 285 926 287
rect 966 285 970 287
rect 860 277 871 279
rect 911 277 926 279
rect 966 277 970 279
rect 285 268 296 270
rect 336 268 351 270
rect 391 268 395 270
rect 285 260 296 262
rect 336 260 351 262
rect 391 260 395 262
rect -37 240 -26 242
rect 14 240 29 242
rect 69 240 73 242
rect 1659 241 1670 243
rect 1710 241 1725 243
rect 1765 241 1769 243
rect -37 232 -26 234
rect 14 232 29 234
rect 69 232 73 234
rect 1659 233 1670 235
rect 1710 233 1725 235
rect 1765 233 1769 235
rect 119 219 130 221
rect 170 219 185 221
rect 225 219 229 221
rect 119 211 130 213
rect 170 211 185 213
rect 225 211 229 213
rect 837 203 848 205
rect 888 203 912 205
rect 992 203 995 205
rect 1825 204 1836 206
rect 1876 204 1891 206
rect 1931 204 1935 206
rect 499 195 501 198
rect 837 195 848 197
rect 888 195 912 197
rect 992 195 995 197
rect 1825 196 1836 198
rect 1876 196 1891 198
rect 1931 196 1935 198
rect 837 187 848 189
rect 888 187 912 189
rect 992 187 995 189
rect 837 179 848 181
rect 888 179 912 181
rect 992 179 995 181
rect 1503 176 1514 178
rect 1554 176 1569 178
rect 1609 176 1613 178
rect 1503 168 1514 170
rect 1554 168 1569 170
rect 1609 168 1613 170
rect 499 141 501 155
rect 1056 154 1067 156
rect 1107 154 1131 156
rect 1211 154 1214 156
rect 1659 155 1670 157
rect 1710 155 1725 157
rect 1765 155 1769 157
rect 1056 146 1067 148
rect 1107 146 1131 148
rect 1211 146 1214 148
rect 1659 147 1670 149
rect 1710 147 1725 149
rect 1765 147 1769 149
rect 91 130 102 132
rect 142 130 157 132
rect 197 130 201 132
rect 91 122 102 124
rect 142 122 157 124
rect 197 122 201 124
rect 1056 138 1067 140
rect 1107 138 1131 140
rect 1211 138 1214 140
rect 1056 130 1067 132
rect 1107 130 1131 132
rect 1211 130 1214 132
rect 499 118 501 121
rect 847 106 858 108
rect 898 106 916 108
rect 976 106 981 108
rect 847 98 858 100
rect 898 98 916 100
rect 976 98 981 100
rect 847 90 858 92
rect 898 90 916 92
rect 976 90 981 92
rect 856 33 867 35
rect 907 33 922 35
rect 962 33 966 35
rect 856 25 867 27
rect 907 25 922 27
rect 962 25 966 27
rect 118 -37 129 -35
rect 169 -37 184 -35
rect 224 -37 228 -35
rect 118 -45 129 -43
rect 169 -45 184 -43
rect 224 -45 228 -43
rect 284 -74 295 -72
rect 335 -74 350 -72
rect 390 -74 394 -72
rect 284 -82 295 -80
rect 335 -82 350 -80
rect 390 -82 394 -80
rect -38 -102 -27 -100
rect 13 -102 28 -100
rect 68 -102 72 -100
rect -38 -110 -27 -108
rect 13 -110 28 -108
rect 68 -110 72 -108
rect 118 -123 129 -121
rect 169 -123 184 -121
rect 224 -123 228 -121
rect 118 -131 129 -129
rect 169 -131 184 -129
rect 224 -131 228 -129
rect 493 -147 495 -144
rect 493 -201 495 -187
rect 90 -212 101 -210
rect 141 -212 156 -210
rect 196 -212 200 -210
rect 90 -220 101 -218
rect 141 -220 156 -218
rect 196 -220 200 -218
rect 493 -224 495 -221
rect 805 -303 816 -301
rect 856 -303 880 -301
rect 960 -303 963 -301
rect 805 -311 816 -309
rect 856 -311 880 -309
rect 960 -311 963 -309
rect 112 -319 123 -317
rect 163 -319 178 -317
rect 218 -319 222 -317
rect 805 -319 816 -317
rect 856 -319 880 -317
rect 960 -319 963 -317
rect 112 -327 123 -325
rect 163 -327 178 -325
rect 218 -327 222 -325
rect 805 -327 816 -325
rect 856 -327 880 -325
rect 960 -327 963 -325
rect 805 -335 816 -333
rect 856 -335 880 -333
rect 960 -335 963 -333
rect 278 -356 289 -354
rect 329 -356 344 -354
rect 384 -356 388 -354
rect 278 -364 289 -362
rect 329 -364 344 -362
rect 384 -364 388 -362
rect -44 -384 -33 -382
rect 7 -384 22 -382
rect 62 -384 66 -382
rect 1089 -388 1100 -386
rect 1140 -388 1164 -386
rect 1244 -388 1247 -386
rect -44 -392 -33 -390
rect 7 -392 22 -390
rect 62 -392 66 -390
rect 1089 -396 1100 -394
rect 1140 -396 1164 -394
rect 1244 -396 1247 -394
rect 112 -405 123 -403
rect 163 -405 178 -403
rect 218 -405 222 -403
rect 1089 -404 1100 -402
rect 1140 -404 1164 -402
rect 1244 -404 1247 -402
rect 112 -413 123 -411
rect 163 -413 178 -411
rect 218 -413 222 -411
rect 1089 -412 1100 -410
rect 1140 -412 1164 -410
rect 1244 -412 1247 -410
rect 1089 -420 1100 -418
rect 1140 -420 1164 -418
rect 1244 -420 1247 -418
rect 827 -464 838 -462
rect 878 -464 902 -462
rect 982 -464 985 -462
rect 827 -472 838 -470
rect 878 -472 902 -470
rect 982 -472 985 -470
rect 827 -480 838 -478
rect 878 -480 902 -478
rect 982 -480 985 -478
rect 827 -488 838 -486
rect 878 -488 902 -486
rect 982 -488 985 -486
rect 84 -494 95 -492
rect 135 -494 150 -492
rect 190 -494 194 -492
rect 84 -502 95 -500
rect 135 -502 150 -500
rect 190 -502 194 -500
rect 840 -608 851 -606
rect 891 -608 909 -606
rect 969 -608 974 -606
rect 840 -616 851 -614
rect 891 -616 909 -614
rect 969 -616 974 -614
rect 840 -624 851 -622
rect 891 -624 909 -622
rect 969 -624 974 -622
rect 860 -698 871 -696
rect 911 -698 926 -696
rect 966 -698 970 -696
rect 860 -706 871 -704
rect 911 -706 926 -704
rect 966 -706 970 -704
<< polycontact >>
rect 138 996 142 1000
rect 138 988 142 992
rect 304 959 308 963
rect 304 951 308 955
rect -18 931 -14 935
rect -18 923 -14 927
rect 138 910 142 914
rect 138 902 142 906
rect 1646 910 1650 914
rect 1646 902 1650 906
rect 1812 873 1816 877
rect 1812 865 1816 869
rect 513 836 517 840
rect 1490 845 1494 849
rect 1490 837 1494 841
rect 110 821 114 825
rect 110 813 114 817
rect 1646 824 1650 828
rect 1646 816 1650 820
rect 145 645 149 649
rect 145 637 149 641
rect 1646 635 1650 639
rect 1646 627 1650 631
rect 311 608 315 612
rect 311 600 315 604
rect 1812 598 1816 602
rect 1812 590 1816 594
rect -11 580 -7 584
rect -11 572 -7 576
rect 853 575 857 579
rect 853 567 857 571
rect 1490 570 1494 574
rect 145 559 149 563
rect 1490 562 1494 566
rect 145 551 149 555
rect 1646 549 1650 553
rect 1646 541 1650 545
rect 1077 510 1081 514
rect 1077 502 1081 506
rect 516 485 520 489
rect 117 470 121 474
rect 117 462 121 466
rect 1648 441 1652 445
rect 1648 433 1652 437
rect 1814 404 1818 408
rect 1814 396 1818 400
rect 1492 376 1496 380
rect 847 368 851 372
rect 847 360 851 364
rect 1492 368 1496 372
rect 847 352 851 356
rect 1648 355 1652 359
rect 1648 347 1652 351
rect 1036 327 1040 331
rect 1036 319 1040 323
rect 115 304 119 308
rect 1036 311 1040 315
rect 115 296 119 300
rect 856 284 860 288
rect 856 276 860 280
rect 281 267 285 271
rect 281 259 285 263
rect -41 239 -37 243
rect 1655 240 1659 244
rect -41 231 -37 235
rect 1655 232 1659 236
rect 115 218 119 222
rect 115 210 119 214
rect 833 202 837 206
rect 1821 203 1825 207
rect 833 194 837 198
rect 1821 195 1825 199
rect 833 186 837 190
rect 833 178 837 182
rect 1499 175 1503 179
rect 1499 167 1503 171
rect 495 144 499 148
rect 1052 153 1056 157
rect 1655 154 1659 158
rect 1052 145 1056 149
rect 1655 146 1659 150
rect 87 129 91 133
rect 87 121 91 125
rect 1052 137 1056 141
rect 1052 129 1056 133
rect 843 105 847 109
rect 843 97 847 101
rect 843 89 847 93
rect 852 32 856 36
rect 852 24 856 28
rect 114 -38 118 -34
rect 114 -46 118 -42
rect 280 -75 284 -71
rect 280 -83 284 -79
rect -42 -103 -38 -99
rect -42 -111 -38 -107
rect 114 -124 118 -120
rect 114 -132 118 -128
rect 489 -198 493 -194
rect 86 -213 90 -209
rect 86 -221 90 -217
rect 801 -304 805 -300
rect 801 -312 805 -308
rect 108 -320 112 -316
rect 108 -328 112 -324
rect 801 -320 805 -316
rect 801 -328 805 -324
rect 801 -336 805 -332
rect 274 -357 278 -353
rect 274 -365 278 -361
rect -48 -385 -44 -381
rect -48 -393 -44 -389
rect 1085 -389 1089 -385
rect 1085 -397 1089 -393
rect 108 -406 112 -402
rect 1085 -405 1089 -401
rect 108 -414 112 -410
rect 1085 -413 1089 -409
rect 1085 -421 1089 -417
rect 823 -465 827 -461
rect 823 -473 827 -469
rect 823 -481 827 -477
rect 80 -495 84 -491
rect 823 -489 827 -485
rect 80 -503 84 -499
rect 836 -609 840 -605
rect 836 -617 840 -613
rect 836 -625 840 -621
rect 856 -699 860 -695
rect 856 -707 860 -703
<< metal1 >>
rect 201 1014 205 1015
rect 201 1010 303 1014
rect 201 1004 205 1010
rect 146 1000 153 1004
rect 201 1000 208 1004
rect 134 999 138 1000
rect -22 996 138 999
rect -22 995 137 996
rect -22 935 -18 995
rect 45 988 138 992
rect 146 988 150 1000
rect 201 996 205 1000
rect 193 992 205 996
rect 45 952 49 988
rect 146 984 153 988
rect 248 984 259 988
rect 141 980 150 984
rect 141 976 145 980
rect 299 963 303 1010
rect 367 977 481 981
rect 367 967 371 977
rect 312 963 319 967
rect 367 963 374 967
rect 299 959 304 963
rect 300 953 304 955
rect 45 948 136 952
rect 45 939 49 948
rect -10 935 -3 939
rect 45 935 52 939
rect -72 931 -51 935
rect -46 931 -18 935
rect -66 923 -18 927
rect -10 923 -6 935
rect 45 931 49 935
rect 37 927 49 931
rect -66 917 -62 923
rect -72 913 -62 917
rect -38 889 -34 923
rect -10 919 -3 923
rect 92 919 103 923
rect -15 915 -6 919
rect -15 911 -11 915
rect 132 914 136 948
rect 201 949 304 953
rect 312 951 316 963
rect 367 959 371 963
rect 359 955 371 959
rect 201 918 205 949
rect 312 947 319 951
rect 414 947 425 951
rect 307 943 316 947
rect 307 939 311 943
rect 1709 928 1713 929
rect 1709 924 1811 928
rect 1709 918 1713 924
rect 146 914 153 918
rect 201 914 208 918
rect 1654 914 1661 918
rect 1709 914 1716 918
rect 132 910 138 914
rect 134 904 138 906
rect 52 902 138 904
rect 146 902 150 914
rect 201 910 205 914
rect 1642 913 1646 914
rect 1486 910 1646 913
rect 193 906 205 910
rect 1486 909 1645 910
rect 52 900 137 902
rect 52 889 56 900
rect -38 885 56 889
rect 97 825 101 900
rect 146 898 153 902
rect 248 898 259 902
rect 141 894 150 898
rect 141 890 145 894
rect 508 893 530 897
rect 512 887 516 893
rect 1486 854 1490 909
rect 1424 850 1490 854
rect 1553 902 1646 906
rect 1654 902 1658 914
rect 1709 910 1713 914
rect 1701 906 1713 910
rect 1553 866 1557 902
rect 1654 898 1661 902
rect 1756 898 1767 902
rect 1649 894 1658 898
rect 1649 890 1653 894
rect 1807 877 1811 924
rect 1875 881 1879 892
rect 1820 877 1827 881
rect 1875 877 1882 881
rect 1807 873 1812 877
rect 1808 867 1812 869
rect 1553 862 1644 866
rect 1553 853 1557 862
rect 520 840 524 847
rect 1486 845 1490 850
rect 1498 849 1505 853
rect 1553 849 1560 853
rect 1465 841 1476 842
rect 173 836 513 840
rect 520 839 538 840
rect 1465 839 1490 841
rect 520 837 1490 839
rect 1498 837 1502 849
rect 1553 845 1557 849
rect 1545 841 1557 845
rect 520 836 1476 837
rect 173 829 177 836
rect 520 833 524 836
rect 118 825 125 829
rect 173 825 180 829
rect 97 821 110 825
rect 109 813 110 817
rect 118 813 122 825
rect 173 821 177 825
rect 165 817 177 821
rect 118 809 125 813
rect 220 809 229 813
rect 534 835 1476 836
rect 113 805 122 809
rect 512 809 516 813
rect 506 805 530 809
rect 113 802 117 805
rect 208 663 212 664
rect 208 659 310 663
rect 208 653 212 659
rect 153 649 160 653
rect 208 649 215 653
rect 141 648 145 649
rect -15 645 145 648
rect -15 644 144 645
rect -15 584 -11 644
rect 52 637 145 641
rect 153 637 157 649
rect 208 645 212 649
rect 200 641 212 645
rect 52 601 56 637
rect 153 633 160 637
rect 255 633 266 637
rect 148 629 157 633
rect 148 625 152 629
rect 306 612 310 659
rect 374 626 498 630
rect 374 616 378 626
rect 319 612 326 616
rect 374 612 381 616
rect 306 608 311 612
rect 307 602 311 604
rect 52 597 143 601
rect 52 588 56 597
rect -3 584 4 588
rect 52 584 59 588
rect -65 580 -44 584
rect -39 580 -11 584
rect -59 572 -11 576
rect -3 572 1 584
rect 52 580 56 584
rect 44 576 56 580
rect -59 566 -55 572
rect -65 562 -55 566
rect -31 538 -27 572
rect -3 568 4 572
rect 99 568 110 572
rect -8 564 1 568
rect -8 560 -4 564
rect 139 563 143 597
rect 208 598 311 602
rect 319 600 323 612
rect 374 608 378 612
rect 366 604 378 608
rect 208 567 212 598
rect 319 596 326 600
rect 421 596 432 600
rect 314 592 323 596
rect 314 588 318 592
rect 484 571 488 626
rect 534 581 538 835
rect 1465 831 1476 835
rect 1498 833 1505 837
rect 1600 833 1611 837
rect 1470 803 1474 831
rect 1493 829 1502 833
rect 1493 825 1497 829
rect 1640 828 1644 862
rect 1709 863 1812 867
rect 1820 865 1824 877
rect 1875 873 1879 877
rect 1867 869 1879 873
rect 1709 832 1713 863
rect 1820 861 1827 865
rect 1922 861 1933 865
rect 1815 857 1824 861
rect 1815 853 1819 857
rect 1654 828 1661 832
rect 1709 828 1716 832
rect 1640 824 1646 828
rect 1642 818 1646 820
rect 1560 816 1646 818
rect 1654 816 1658 828
rect 1709 824 1713 828
rect 1701 820 1713 824
rect 1560 814 1645 816
rect 1560 803 1564 814
rect 1654 812 1661 816
rect 1756 812 1767 816
rect 1649 808 1658 812
rect 1649 804 1653 808
rect 1470 799 1564 803
rect 1709 653 1713 654
rect 1709 649 1811 653
rect 1709 643 1713 649
rect 1654 639 1661 643
rect 1709 639 1716 643
rect 1642 638 1646 639
rect 1486 635 1646 638
rect 1486 634 1645 635
rect 672 581 676 584
rect 916 586 1040 590
rect 916 583 920 586
rect 534 579 852 581
rect 861 579 868 583
rect 916 579 923 583
rect 534 577 820 579
rect 825 577 853 579
rect 843 575 853 577
rect 843 574 852 575
rect 484 567 853 571
rect 861 567 865 579
rect 916 575 920 579
rect 908 571 920 575
rect 153 563 160 567
rect 208 563 215 567
rect 747 564 751 567
rect 829 564 833 567
rect 139 559 145 563
rect 141 553 145 555
rect 59 551 145 553
rect 153 551 157 563
rect 208 559 212 563
rect 861 563 868 567
rect 963 563 972 567
rect 856 559 865 563
rect 200 555 212 559
rect 856 556 860 559
rect 59 549 144 551
rect 59 538 63 549
rect -31 534 63 538
rect 104 474 108 549
rect 153 547 160 551
rect 255 547 266 551
rect 148 543 157 547
rect 148 539 152 543
rect 511 542 533 546
rect 515 536 519 542
rect 1036 514 1040 586
rect 1486 574 1490 634
rect 1553 627 1646 631
rect 1654 627 1658 639
rect 1709 635 1713 639
rect 1701 631 1713 635
rect 1553 591 1557 627
rect 1654 623 1661 627
rect 1756 623 1767 627
rect 1649 619 1658 623
rect 1649 615 1653 619
rect 1807 602 1811 649
rect 1875 606 1879 617
rect 1820 602 1827 606
rect 1875 602 1882 606
rect 1807 598 1812 602
rect 1808 592 1812 594
rect 1553 587 1644 591
rect 1553 578 1557 587
rect 1498 574 1505 578
rect 1553 574 1560 578
rect 1437 570 1490 574
rect 1437 569 1489 570
rect 1470 565 1490 566
rect 1384 562 1490 565
rect 1498 562 1502 574
rect 1553 570 1557 574
rect 1545 566 1557 570
rect 1384 561 1475 562
rect 1384 542 1388 561
rect 1140 538 1388 542
rect 1140 518 1144 538
rect 1085 514 1092 518
rect 1140 514 1147 518
rect 1036 510 1077 514
rect 523 489 527 496
rect 1036 502 1077 506
rect 1085 502 1089 514
rect 1140 510 1144 514
rect 1132 506 1144 510
rect 180 485 516 489
rect 523 487 811 489
rect 523 485 759 487
rect 180 478 184 485
rect 125 474 132 478
rect 180 474 187 478
rect 104 470 117 474
rect 116 462 117 466
rect 125 462 129 474
rect 180 470 184 474
rect 172 466 184 470
rect 125 458 132 462
rect 227 458 236 462
rect 120 454 129 458
rect 120 451 124 454
rect 461 442 465 485
rect 523 482 527 485
rect 581 478 585 485
rect 764 485 811 487
rect 515 458 519 462
rect 509 454 533 458
rect 553 446 898 450
rect 1036 442 1040 502
rect 1085 498 1092 502
rect 1187 498 1196 502
rect 1080 494 1089 498
rect 1080 491 1084 494
rect 461 438 1040 442
rect 178 322 182 323
rect 178 318 280 322
rect 178 312 182 318
rect 123 308 130 312
rect 178 308 185 312
rect 111 307 115 308
rect -45 304 115 307
rect -45 303 114 304
rect -45 243 -41 303
rect 22 296 115 300
rect 123 296 127 308
rect 178 304 182 308
rect 170 300 182 304
rect 22 260 26 296
rect 123 292 130 296
rect 225 292 236 296
rect 118 288 127 292
rect 118 284 122 288
rect 276 271 280 318
rect 548 289 552 420
rect 820 364 824 423
rect 829 372 833 423
rect 898 420 902 424
rect 1432 420 1436 543
rect 1470 528 1474 561
rect 1498 558 1505 562
rect 1600 558 1611 562
rect 1493 554 1502 558
rect 1493 550 1497 554
rect 1640 553 1644 587
rect 1709 588 1812 592
rect 1820 590 1824 602
rect 1875 598 1879 602
rect 1867 594 1879 598
rect 1709 557 1713 588
rect 1820 586 1827 590
rect 1922 586 1933 590
rect 1815 582 1824 586
rect 1815 578 1819 582
rect 1654 553 1661 557
rect 1709 553 1716 557
rect 1640 549 1646 553
rect 1642 543 1646 545
rect 1560 541 1646 543
rect 1654 541 1658 553
rect 1709 549 1713 553
rect 1701 545 1713 549
rect 1560 539 1645 541
rect 1560 528 1564 539
rect 1654 537 1661 541
rect 1756 537 1767 541
rect 1649 533 1658 537
rect 1649 529 1653 533
rect 1470 524 1564 528
rect 1711 459 1715 460
rect 1711 455 1813 459
rect 1711 449 1715 455
rect 1656 445 1663 449
rect 1711 445 1718 449
rect 1644 444 1648 445
rect 898 416 1436 420
rect 1488 441 1648 444
rect 1488 440 1647 441
rect 1104 379 1390 383
rect 902 372 920 376
rect 829 368 847 372
rect 855 364 862 368
rect 820 360 847 364
rect 796 352 847 356
rect 855 352 859 364
rect 906 360 910 372
rect 902 356 910 360
rect 796 289 800 352
rect 855 348 862 352
rect 855 342 859 348
rect 906 331 910 356
rect 980 348 997 352
rect 1104 335 1108 379
rect 1386 372 1390 379
rect 1488 382 1492 440
rect 1555 433 1648 437
rect 1656 433 1660 445
rect 1711 441 1715 445
rect 1703 437 1715 441
rect 1555 397 1559 433
rect 1656 429 1663 433
rect 1758 429 1769 433
rect 1651 425 1660 429
rect 1651 421 1655 425
rect 1809 408 1813 455
rect 1877 412 1881 423
rect 1822 408 1829 412
rect 1877 408 1884 412
rect 1809 404 1814 408
rect 1810 398 1814 400
rect 1555 393 1646 397
rect 1555 384 1559 393
rect 1456 378 1492 382
rect 1500 380 1507 384
rect 1555 380 1562 384
rect 1488 376 1492 378
rect 1386 368 1492 372
rect 1500 368 1504 380
rect 1555 376 1559 380
rect 1547 372 1559 376
rect 1091 331 1109 335
rect 1472 334 1476 368
rect 1500 364 1507 368
rect 1602 364 1613 368
rect 1495 360 1504 364
rect 1495 356 1499 360
rect 1642 359 1646 393
rect 1711 394 1814 398
rect 1822 396 1826 408
rect 1877 404 1881 408
rect 1869 400 1881 404
rect 1711 363 1715 394
rect 1822 392 1829 396
rect 1924 392 1935 396
rect 1817 388 1826 392
rect 1817 384 1821 388
rect 1656 359 1663 363
rect 1711 359 1718 363
rect 1642 355 1648 359
rect 1644 349 1648 351
rect 1562 347 1648 349
rect 1656 347 1660 359
rect 1711 355 1715 359
rect 1703 351 1715 355
rect 1562 345 1647 347
rect 1562 334 1566 345
rect 1656 343 1663 347
rect 1758 343 1769 347
rect 1651 339 1660 343
rect 1651 335 1655 339
rect 906 327 1036 331
rect 1044 323 1051 327
rect 919 319 1036 323
rect 919 292 923 319
rect 1000 311 1036 315
rect 1044 311 1048 323
rect 1095 319 1099 331
rect 1472 330 1566 334
rect 1091 315 1099 319
rect 1044 307 1051 311
rect 1169 307 1186 311
rect 1044 301 1048 307
rect 344 288 842 289
rect 864 288 871 292
rect 919 288 926 292
rect 344 285 856 288
rect 344 275 348 285
rect 622 284 631 285
rect 627 283 631 284
rect 289 271 296 275
rect 344 271 351 275
rect 467 271 794 275
rect 276 267 281 271
rect 277 261 281 263
rect 22 256 113 260
rect 22 247 26 256
rect -33 243 -26 247
rect 22 243 29 247
rect -95 239 -74 243
rect -69 239 -41 243
rect -89 231 -41 235
rect -33 231 -29 243
rect 22 239 26 243
rect 14 235 26 239
rect -89 225 -85 231
rect -95 221 -85 225
rect -61 197 -57 231
rect -33 227 -26 231
rect 69 227 80 231
rect -38 223 -29 227
rect -38 219 -34 223
rect 109 222 113 256
rect 178 257 281 261
rect 289 259 293 271
rect 344 267 348 271
rect 336 263 348 267
rect 178 226 182 257
rect 289 255 296 259
rect 391 255 402 259
rect 284 251 293 255
rect 284 247 288 251
rect 123 222 130 226
rect 178 222 185 226
rect 109 218 115 222
rect 111 212 115 214
rect 29 210 115 212
rect 123 210 127 222
rect 178 218 182 222
rect 170 214 182 218
rect 29 208 114 210
rect 29 197 33 208
rect -61 193 33 197
rect 74 133 78 208
rect 123 206 130 210
rect 225 206 236 210
rect 118 202 127 206
rect 118 198 122 202
rect 467 148 471 271
rect 747 206 751 255
rect 802 215 806 285
rect 838 284 856 285
rect 816 276 856 280
rect 864 276 868 288
rect 919 284 923 288
rect 911 280 923 284
rect 864 272 871 276
rect 966 272 975 276
rect 859 268 868 272
rect 859 265 863 268
rect 1718 258 1722 259
rect 1718 254 1820 258
rect 1718 248 1722 254
rect 1663 244 1670 248
rect 1718 244 1725 248
rect 1651 243 1655 244
rect 1495 240 1655 243
rect 1495 239 1654 240
rect 840 206 848 210
rect 891 206 912 210
rect 492 201 512 205
rect 747 202 833 206
rect 494 195 498 201
rect 782 194 833 198
rect 840 194 845 206
rect 891 202 895 206
rect 888 198 895 202
rect 840 190 848 194
rect 807 186 833 190
rect 828 181 833 182
rect 502 148 506 155
rect 797 178 833 181
rect 840 178 845 190
rect 891 186 895 198
rect 1118 193 1394 197
rect 888 182 895 186
rect 797 177 832 178
rect 150 144 495 148
rect 502 144 744 148
rect 150 137 154 144
rect 502 141 506 144
rect 95 133 102 137
rect 150 133 157 137
rect 74 129 87 133
rect 86 121 87 125
rect 95 121 99 133
rect 150 129 154 133
rect 142 125 154 129
rect 95 117 102 121
rect 197 117 206 121
rect 568 139 572 144
rect 90 113 99 117
rect 494 117 498 121
rect 491 113 512 117
rect 90 110 94 113
rect 740 108 744 144
rect 797 94 801 177
rect 840 174 848 178
rect 840 164 845 174
rect 891 167 895 182
rect 992 174 1013 178
rect 891 163 1047 167
rect 1043 157 1047 163
rect 1118 161 1122 193
rect 1390 171 1394 193
rect 1495 181 1499 239
rect 1562 232 1655 236
rect 1663 232 1667 244
rect 1718 240 1722 244
rect 1710 236 1722 240
rect 1562 196 1566 232
rect 1663 228 1670 232
rect 1765 228 1776 232
rect 1658 224 1667 228
rect 1658 220 1662 224
rect 1816 207 1820 254
rect 1884 211 1888 222
rect 1829 207 1836 211
rect 1884 207 1891 211
rect 1816 203 1821 207
rect 1817 197 1821 199
rect 1562 192 1653 196
rect 1562 183 1566 192
rect 1447 177 1499 181
rect 1507 179 1514 183
rect 1562 179 1569 183
rect 1495 175 1499 177
rect 1390 167 1499 171
rect 1507 167 1511 179
rect 1562 175 1566 179
rect 1554 171 1566 175
rect 1059 157 1067 161
rect 1110 157 1131 161
rect 1043 153 1052 157
rect 907 145 1052 149
rect 1059 145 1064 157
rect 1110 153 1114 157
rect 1107 149 1114 153
rect 907 113 911 145
rect 1059 141 1067 145
rect 1027 137 1052 141
rect 898 109 916 113
rect 836 105 843 109
rect 851 101 858 105
rect 826 97 843 101
rect 453 93 839 94
rect 453 90 843 93
rect 453 2 457 90
rect 548 85 552 90
rect 740 29 744 82
rect 816 37 820 90
rect 835 89 843 90
rect 851 89 855 101
rect 902 97 906 109
rect 898 93 906 97
rect 851 85 858 89
rect 976 85 993 89
rect 851 79 855 85
rect 1027 62 1031 137
rect 915 58 1031 62
rect 1043 129 1052 133
rect 1059 129 1064 141
rect 1110 137 1114 149
rect 1107 133 1114 137
rect 915 40 919 58
rect 816 36 846 37
rect 860 36 867 40
rect 915 36 922 40
rect 816 33 852 36
rect 842 32 852 33
rect 740 28 848 29
rect 740 25 852 28
rect 842 24 852 25
rect 860 24 864 36
rect 915 32 919 36
rect 907 28 919 32
rect 860 20 867 24
rect 962 20 971 24
rect 855 16 864 20
rect 855 13 859 16
rect 1043 12 1047 129
rect 1059 125 1067 129
rect 1211 125 1229 129
rect 1062 119 1066 125
rect 453 -2 1020 2
rect 177 -20 181 -19
rect 177 -24 279 -20
rect 177 -30 181 -24
rect 122 -34 129 -30
rect 177 -34 184 -30
rect 110 -35 114 -34
rect -46 -38 114 -35
rect -46 -39 113 -38
rect -46 -99 -42 -39
rect 21 -46 114 -42
rect 122 -46 126 -34
rect 177 -38 181 -34
rect 169 -42 181 -38
rect 21 -82 25 -46
rect 122 -50 129 -46
rect 224 -50 235 -46
rect 117 -54 126 -50
rect 117 -58 121 -54
rect 275 -71 279 -24
rect 453 -53 457 -2
rect 1041 -5 1047 12
rect 1041 -18 1045 -5
rect 343 -57 457 -53
rect 487 -22 1045 -18
rect 343 -67 347 -57
rect 288 -71 295 -67
rect 343 -71 350 -67
rect 275 -75 280 -71
rect 276 -81 280 -79
rect 21 -86 112 -82
rect 21 -95 25 -86
rect -34 -99 -27 -95
rect 21 -99 28 -95
rect -96 -103 -75 -99
rect -70 -103 -42 -99
rect -90 -111 -42 -107
rect -34 -111 -30 -99
rect 21 -103 25 -99
rect 13 -107 25 -103
rect -90 -117 -86 -111
rect -96 -121 -86 -117
rect -62 -145 -58 -111
rect -34 -115 -27 -111
rect 68 -115 79 -111
rect -39 -119 -30 -115
rect -39 -123 -35 -119
rect 108 -120 112 -86
rect 177 -85 280 -81
rect 288 -83 292 -71
rect 343 -75 347 -71
rect 335 -79 347 -75
rect 487 -78 491 -22
rect 454 -82 491 -78
rect 177 -116 181 -85
rect 288 -87 295 -83
rect 390 -87 401 -83
rect 283 -91 292 -87
rect 283 -95 287 -91
rect 122 -120 129 -116
rect 177 -120 184 -116
rect 108 -124 114 -120
rect 110 -130 114 -128
rect 28 -132 114 -130
rect 122 -132 126 -120
rect 177 -124 181 -120
rect 169 -128 181 -124
rect 28 -134 113 -132
rect 28 -145 32 -134
rect -62 -149 32 -145
rect 73 -209 77 -134
rect 122 -136 129 -132
rect 224 -136 235 -132
rect 117 -140 126 -136
rect 117 -144 121 -140
rect 454 -194 458 -82
rect 483 -141 506 -137
rect 488 -147 492 -141
rect 496 -194 500 -187
rect 149 -198 489 -194
rect 496 -198 514 -194
rect 149 -205 153 -198
rect 496 -201 500 -198
rect 94 -209 101 -205
rect 149 -209 156 -205
rect 73 -213 86 -209
rect 85 -221 86 -217
rect 94 -221 98 -209
rect 149 -213 153 -209
rect 141 -217 153 -213
rect 94 -225 101 -221
rect 196 -225 205 -221
rect 89 -229 98 -225
rect 488 -225 492 -221
rect 482 -229 506 -225
rect 89 -232 93 -229
rect 171 -302 175 -301
rect 171 -306 273 -302
rect 171 -312 175 -306
rect 116 -316 123 -312
rect 171 -316 178 -312
rect 104 -317 108 -316
rect -52 -320 108 -317
rect -52 -321 107 -320
rect -52 -381 -48 -321
rect 15 -328 108 -324
rect 116 -328 120 -316
rect 171 -320 175 -316
rect 163 -324 175 -320
rect 15 -364 19 -328
rect 116 -332 123 -328
rect 218 -332 229 -328
rect 111 -336 120 -332
rect 111 -340 115 -336
rect 269 -353 273 -306
rect 510 -322 514 -198
rect 1442 -202 1446 150
rect 1479 133 1483 167
rect 1507 163 1514 167
rect 1609 163 1620 167
rect 1502 159 1511 163
rect 1502 155 1506 159
rect 1649 158 1653 192
rect 1718 193 1821 197
rect 1829 195 1833 207
rect 1884 203 1888 207
rect 1876 199 1888 203
rect 1718 162 1722 193
rect 1829 191 1836 195
rect 1931 191 1942 195
rect 1824 187 1833 191
rect 1824 183 1828 187
rect 1663 158 1670 162
rect 1718 158 1725 162
rect 1649 154 1655 158
rect 1651 148 1655 150
rect 1569 146 1655 148
rect 1663 146 1667 158
rect 1718 154 1722 158
rect 1710 150 1722 154
rect 1569 144 1654 146
rect 1569 133 1573 144
rect 1663 142 1670 146
rect 1765 142 1776 146
rect 1658 138 1667 142
rect 1658 134 1662 138
rect 1479 129 1573 133
rect 529 -206 1446 -202
rect 529 -335 533 -206
rect 658 -285 800 -281
rect 796 -300 800 -285
rect 856 -300 880 -296
rect 796 -304 801 -300
rect 808 -308 816 -304
rect 712 -312 801 -308
rect 662 -320 801 -316
rect 808 -320 812 -308
rect 861 -312 865 -300
rect 856 -316 865 -312
rect 808 -324 816 -320
rect 561 -328 801 -324
rect 770 -335 801 -332
rect 337 -336 801 -335
rect 808 -336 812 -324
rect 861 -328 865 -316
rect 856 -332 865 -328
rect 337 -339 774 -336
rect 337 -349 341 -339
rect 282 -353 289 -349
rect 337 -353 344 -349
rect 447 -350 451 -339
rect 808 -340 816 -336
rect 808 -349 812 -340
rect 269 -357 274 -353
rect 270 -363 274 -361
rect 15 -368 106 -364
rect 15 -377 19 -368
rect -40 -381 -33 -377
rect 15 -381 22 -377
rect -102 -385 -81 -381
rect -76 -385 -48 -381
rect -96 -393 -48 -389
rect -40 -393 -36 -381
rect 15 -385 19 -381
rect 7 -389 19 -385
rect -96 -399 -92 -393
rect -102 -403 -92 -399
rect -68 -427 -64 -393
rect -40 -397 -33 -393
rect 62 -397 73 -393
rect -45 -401 -36 -397
rect -45 -405 -41 -401
rect 102 -402 106 -368
rect 171 -367 274 -363
rect 282 -365 286 -353
rect 337 -357 341 -353
rect 868 -353 872 -300
rect 960 -340 980 -336
rect 868 -357 1084 -353
rect 329 -361 341 -357
rect 171 -398 175 -367
rect 282 -369 289 -365
rect 384 -369 395 -365
rect 277 -373 286 -369
rect 277 -377 281 -373
rect 510 -390 514 -357
rect 936 -380 1063 -376
rect 1059 -393 1063 -380
rect 1080 -385 1084 -357
rect 1153 -361 1490 -357
rect 1153 -381 1157 -361
rect 1140 -385 1164 -381
rect 1080 -389 1085 -385
rect 1092 -393 1100 -389
rect 1059 -397 1085 -393
rect 116 -402 123 -398
rect 171 -402 178 -398
rect 863 -401 1033 -397
rect 102 -406 108 -402
rect 104 -412 108 -410
rect 22 -414 108 -412
rect 116 -414 120 -402
rect 171 -406 175 -402
rect 163 -410 175 -406
rect 863 -410 867 -401
rect 1029 -402 1033 -401
rect 1080 -402 1085 -401
rect 1029 -406 1085 -402
rect 1092 -405 1096 -393
rect 1145 -397 1149 -385
rect 1140 -401 1149 -397
rect 1092 -409 1100 -405
rect 22 -416 107 -414
rect 22 -427 26 -416
rect -68 -431 26 -427
rect 67 -491 71 -416
rect 116 -418 123 -414
rect 218 -418 229 -414
rect 449 -414 867 -410
rect 907 -413 1085 -409
rect 111 -422 120 -418
rect 111 -426 115 -422
rect 449 -476 453 -414
rect 890 -421 1085 -417
rect 1092 -421 1096 -409
rect 1145 -413 1149 -401
rect 1140 -417 1149 -413
rect 143 -480 453 -476
rect 143 -487 147 -480
rect 88 -491 95 -487
rect 143 -491 150 -487
rect 67 -495 80 -491
rect 79 -503 80 -499
rect 88 -503 92 -491
rect 143 -495 147 -491
rect 135 -499 147 -495
rect 88 -507 95 -503
rect 190 -507 199 -503
rect 83 -511 92 -507
rect 83 -514 87 -511
rect 510 -666 514 -433
rect 600 -458 822 -454
rect 890 -457 894 -421
rect 1092 -425 1100 -421
rect 1244 -425 1264 -421
rect 1092 -434 1096 -425
rect 818 -461 822 -458
rect 830 -461 838 -457
rect 881 -461 902 -457
rect 818 -465 823 -461
rect 713 -473 823 -469
rect 830 -473 835 -461
rect 881 -465 885 -461
rect 878 -469 885 -465
rect 830 -477 838 -473
rect 754 -481 823 -477
rect 754 -617 758 -481
rect 802 -489 823 -485
rect 830 -489 835 -477
rect 881 -481 885 -469
rect 878 -485 885 -481
rect 802 -620 806 -489
rect 830 -493 838 -489
rect 982 -493 1000 -489
rect 833 -499 837 -493
rect 900 -601 904 -587
rect 891 -605 909 -601
rect 830 -609 836 -605
rect 844 -613 851 -609
rect 819 -617 836 -613
rect 802 -621 832 -620
rect 802 -624 836 -621
rect 510 -670 770 -666
rect 802 -703 806 -624
rect 829 -625 836 -624
rect 844 -625 848 -613
rect 895 -617 899 -605
rect 891 -621 899 -617
rect 844 -629 851 -625
rect 969 -629 986 -625
rect 844 -635 848 -629
rect 833 -695 837 -671
rect 919 -691 923 -676
rect 864 -695 871 -691
rect 919 -695 926 -691
rect 833 -699 856 -695
rect 792 -707 856 -703
rect 864 -707 868 -695
rect 919 -699 923 -695
rect 911 -703 923 -699
rect 864 -711 871 -707
rect 966 -711 975 -707
rect 859 -715 868 -711
rect 859 -718 863 -715
<< m2contact >>
rect 259 984 264 989
rect 140 971 145 976
rect -51 930 -46 935
rect 103 919 108 924
rect -16 906 -11 911
rect 425 947 430 952
rect 306 934 311 939
rect 259 898 264 903
rect 503 893 508 898
rect 140 885 145 890
rect 1418 850 1424 856
rect 1767 898 1772 903
rect 1648 885 1653 890
rect 104 812 109 817
rect 229 809 234 814
rect 501 805 506 810
rect 112 797 117 802
rect 266 633 271 638
rect 147 620 152 625
rect 498 626 503 631
rect -44 579 -39 584
rect 110 568 115 573
rect -9 555 -4 560
rect 432 596 437 601
rect 313 583 318 588
rect 1611 833 1616 838
rect 1492 820 1497 825
rect 1933 861 1938 866
rect 1814 848 1819 853
rect 1767 812 1772 817
rect 1648 799 1653 804
rect 671 584 676 589
rect 820 574 825 579
rect 747 559 752 564
rect 829 559 834 564
rect 972 563 977 568
rect 266 547 271 552
rect 855 551 860 556
rect 506 542 511 547
rect 147 534 152 539
rect 1767 623 1772 628
rect 1648 610 1653 615
rect 1432 569 1437 574
rect 1432 543 1437 548
rect 111 461 116 466
rect 236 458 241 463
rect 119 446 124 451
rect 759 482 764 487
rect 811 485 816 490
rect 581 473 586 478
rect 504 454 509 459
rect 548 446 553 451
rect 898 446 903 451
rect 1196 498 1201 503
rect 1079 486 1084 491
rect 548 420 553 425
rect 820 423 825 428
rect 829 423 834 428
rect 898 424 903 429
rect 236 292 241 297
rect 117 279 122 284
rect 1611 558 1616 563
rect 1492 545 1497 550
rect 1933 586 1938 591
rect 1814 573 1819 578
rect 1767 537 1772 542
rect 1648 524 1653 529
rect 854 337 859 342
rect 997 348 1002 353
rect 1451 378 1456 383
rect 1769 429 1774 434
rect 1650 416 1655 421
rect 1613 364 1618 369
rect 1494 351 1499 356
rect 1935 392 1940 397
rect 1816 379 1821 384
rect 1769 343 1774 348
rect 995 311 1000 316
rect 1650 330 1655 335
rect 1186 307 1191 312
rect 1043 296 1048 301
rect 622 279 627 284
rect 794 271 799 276
rect -74 238 -69 243
rect 80 227 85 232
rect -39 214 -34 219
rect 402 255 407 260
rect 283 242 288 247
rect 236 206 241 211
rect 117 193 122 198
rect 747 255 752 260
rect 811 276 816 281
rect 975 272 980 277
rect 858 260 863 265
rect 802 210 807 215
rect 487 201 492 206
rect 777 193 782 198
rect 802 185 807 190
rect 81 120 86 125
rect 206 117 211 122
rect 568 134 573 139
rect 486 113 491 118
rect 89 105 94 110
rect 740 103 745 108
rect 840 159 845 164
rect 1013 174 1018 179
rect 1776 228 1781 233
rect 1657 215 1662 220
rect 1442 176 1447 181
rect 1442 150 1447 155
rect 831 105 836 110
rect 821 97 826 102
rect 548 80 553 85
rect 740 82 745 87
rect 993 85 998 90
rect 850 74 855 79
rect 971 20 976 25
rect 854 8 859 13
rect 1229 125 1234 130
rect 1061 114 1066 119
rect 1020 -2 1025 3
rect 235 -50 240 -45
rect 116 -63 121 -58
rect -75 -104 -70 -99
rect 79 -115 84 -110
rect -40 -128 -35 -123
rect 401 -87 406 -82
rect 282 -100 287 -95
rect 235 -136 240 -131
rect 116 -149 121 -144
rect 478 -141 483 -136
rect 80 -222 85 -217
rect 205 -225 210 -220
rect 477 -229 482 -224
rect 88 -237 93 -232
rect 229 -332 234 -327
rect 110 -345 115 -340
rect 1620 163 1625 168
rect 1501 150 1506 155
rect 1942 191 1947 196
rect 1823 178 1828 183
rect 1776 142 1781 147
rect 1657 129 1662 134
rect 510 -327 515 -322
rect 653 -285 658 -280
rect 712 -308 717 -303
rect 657 -320 662 -315
rect 556 -328 561 -323
rect -81 -386 -76 -381
rect 73 -397 78 -392
rect -46 -410 -41 -405
rect 447 -355 452 -350
rect 510 -357 515 -352
rect 807 -354 812 -349
rect 980 -340 985 -335
rect 395 -369 400 -364
rect 276 -382 281 -377
rect 931 -380 936 -375
rect 510 -395 515 -390
rect 229 -418 234 -413
rect 902 -414 907 -409
rect 110 -431 115 -426
rect 510 -433 515 -428
rect 74 -504 79 -499
rect 199 -507 204 -502
rect 82 -519 87 -514
rect 595 -458 600 -453
rect 1264 -425 1269 -420
rect 1091 -439 1096 -434
rect 708 -473 713 -467
rect 754 -622 759 -617
rect 1000 -493 1005 -488
rect 832 -504 837 -499
rect 900 -587 905 -582
rect 825 -609 830 -604
rect 814 -617 819 -612
rect 770 -670 775 -665
rect 786 -707 792 -701
rect 986 -629 991 -624
rect 843 -640 848 -635
rect 833 -671 838 -666
rect 919 -676 924 -671
rect 975 -711 980 -706
rect 858 -723 863 -718
<< metal2 >>
rect 260 989 264 993
rect 135 971 140 975
rect 426 952 430 956
rect 301 934 306 938
rect -51 817 -47 930
rect 104 924 108 928
rect -21 906 -16 910
rect 260 903 264 907
rect 1768 903 1772 907
rect 499 893 503 897
rect 135 885 140 889
rect 1643 885 1648 889
rect 1934 866 1938 870
rect 1224 850 1418 854
rect -51 813 104 817
rect 230 814 234 818
rect 497 805 501 809
rect 108 797 112 801
rect 267 638 271 642
rect 1224 630 1228 850
rect 1809 848 1814 852
rect 1612 838 1616 842
rect 1487 820 1492 824
rect 1768 817 1772 821
rect 1643 799 1648 803
rect 503 626 1228 630
rect 1768 628 1772 632
rect 142 620 147 624
rect 1643 610 1648 614
rect 433 601 437 605
rect 643 602 676 606
rect 308 583 313 587
rect -44 466 -40 579
rect 111 573 115 577
rect -14 555 -9 559
rect 267 552 271 556
rect 502 542 506 546
rect 142 534 147 538
rect -44 462 111 466
rect 237 463 241 467
rect 500 454 504 458
rect 115 446 119 450
rect 548 425 552 446
rect 237 297 241 301
rect 112 279 117 283
rect 403 260 407 264
rect 278 242 283 246
rect -74 125 -70 238
rect 81 232 85 236
rect -44 214 -39 218
rect 237 211 241 215
rect 483 201 487 205
rect 112 193 117 197
rect -74 121 81 125
rect 207 122 211 126
rect 482 113 486 117
rect 85 105 89 109
rect 236 -45 240 -41
rect 111 -63 116 -59
rect 402 -82 406 -78
rect 277 -100 282 -96
rect -75 -217 -71 -104
rect 80 -110 84 -106
rect -45 -128 -40 -124
rect 236 -131 240 -127
rect 474 -141 478 -137
rect 111 -149 116 -145
rect -75 -221 80 -217
rect 206 -220 210 -216
rect 473 -229 477 -225
rect 84 -237 88 -233
rect 230 -327 234 -323
rect 548 -324 552 80
rect 105 -345 110 -341
rect 510 -352 514 -327
rect 548 -328 556 -324
rect 396 -364 400 -360
rect 271 -382 276 -378
rect -81 -499 -77 -386
rect 74 -392 78 -388
rect -51 -410 -46 -406
rect 230 -413 234 -409
rect 105 -431 110 -427
rect -81 -503 74 -499
rect 200 -502 204 -498
rect 78 -519 82 -515
rect 447 -705 451 -355
rect 510 -428 514 -395
rect 548 -625 552 -328
rect 568 -602 572 134
rect 581 -454 585 473
rect 622 -316 626 279
rect 643 -281 647 602
rect 672 589 676 602
rect 1934 591 1938 595
rect 747 349 751 559
rect 820 531 824 574
rect 973 568 977 572
rect 777 527 824 531
rect 679 345 751 349
rect 643 -285 653 -281
rect 679 -303 683 345
rect 747 260 751 345
rect 740 87 744 103
rect 759 101 763 482
rect 777 198 781 527
rect 811 281 815 485
rect 820 428 824 527
rect 1809 573 1814 577
rect 829 428 833 559
rect 851 551 855 555
rect 1432 548 1436 569
rect 1612 563 1616 567
rect 1487 545 1492 549
rect 1768 542 1772 546
rect 1643 524 1648 528
rect 1197 503 1201 507
rect 1075 486 1079 490
rect 898 429 902 446
rect 1770 434 1774 438
rect 1645 416 1650 420
rect 1936 397 1940 401
rect 1285 393 1439 397
rect 998 353 1002 357
rect 850 337 854 341
rect 820 311 995 315
rect 1187 312 1191 316
rect 820 272 823 311
rect 1039 296 1043 300
rect 976 277 980 281
rect 799 271 823 272
rect 794 268 823 271
rect 854 260 858 264
rect 802 190 806 210
rect 802 109 806 185
rect 1014 179 1018 183
rect 836 159 840 163
rect 1230 130 1234 134
rect 1057 114 1061 118
rect 802 106 831 109
rect 802 105 817 106
rect 830 105 831 106
rect 759 97 821 101
rect 994 90 998 94
rect 846 74 850 78
rect 972 25 976 29
rect 850 8 854 12
rect 1285 2 1289 393
rect 1435 382 1439 393
rect 1435 378 1451 382
rect 1811 379 1816 383
rect 1614 369 1618 373
rect 1489 351 1494 355
rect 1770 348 1774 352
rect 1645 330 1650 334
rect 1777 233 1781 237
rect 1652 215 1657 219
rect 1943 196 1947 200
rect 1818 178 1823 182
rect 1442 155 1446 176
rect 1621 168 1625 172
rect 1496 150 1501 154
rect 1777 147 1781 151
rect 1652 129 1657 133
rect 1025 -2 1289 2
rect 679 -307 712 -303
rect 622 -320 657 -316
rect 581 -458 595 -454
rect 622 -471 626 -320
rect 981 -335 985 -331
rect 803 -354 807 -350
rect 919 -380 931 -376
rect 900 -414 902 -409
rect 693 -471 708 -467
rect 622 -475 697 -471
rect 828 -504 832 -500
rect 900 -582 904 -414
rect 568 -604 830 -602
rect 568 -606 825 -604
rect 768 -617 814 -613
rect 768 -621 772 -617
rect 759 -622 772 -621
rect 754 -625 772 -622
rect 548 -629 772 -625
rect 839 -640 843 -636
rect 775 -670 833 -666
rect 919 -671 923 -380
rect 1265 -420 1269 -416
rect 1087 -439 1091 -435
rect 1001 -488 1005 -484
rect 987 -624 991 -620
rect 447 -707 786 -705
rect 976 -706 980 -702
rect 447 -709 790 -707
rect 854 -723 858 -719
<< m3contact >>
rect 259 993 264 998
rect 130 971 135 976
rect 425 956 430 961
rect 296 934 301 939
rect 103 928 108 933
rect -26 906 -21 911
rect 259 907 264 912
rect 1767 907 1772 912
rect 494 893 499 898
rect 130 885 135 890
rect 1638 885 1643 890
rect 1933 870 1938 875
rect 229 818 234 823
rect 492 805 497 810
rect 103 797 108 802
rect 266 642 271 647
rect 1804 848 1809 853
rect 1611 842 1616 847
rect 1482 820 1487 825
rect 1767 821 1772 826
rect 1638 799 1643 804
rect 1767 632 1772 637
rect 137 620 142 625
rect 1638 610 1643 615
rect 432 605 437 610
rect 303 583 308 588
rect 110 577 115 582
rect -19 555 -14 560
rect 266 556 271 561
rect 497 542 502 547
rect 137 534 142 539
rect 236 467 241 472
rect 495 454 500 459
rect 110 446 115 451
rect 236 301 241 306
rect 107 279 112 284
rect 402 264 407 269
rect 273 242 278 247
rect 80 236 85 241
rect -49 214 -44 219
rect 236 215 241 220
rect 478 201 483 206
rect 107 193 112 198
rect 206 126 211 131
rect 477 113 482 118
rect 80 105 85 110
rect 235 -41 240 -36
rect 106 -63 111 -58
rect 401 -78 406 -73
rect 272 -100 277 -95
rect 79 -106 84 -101
rect -50 -128 -45 -123
rect 235 -127 240 -122
rect 469 -141 474 -136
rect 106 -149 111 -144
rect 205 -216 210 -211
rect 468 -229 473 -224
rect 79 -237 84 -232
rect 229 -323 234 -318
rect 100 -345 105 -340
rect 395 -360 400 -355
rect 266 -382 271 -377
rect 73 -388 78 -383
rect -56 -410 -51 -405
rect 229 -409 234 -404
rect 100 -431 105 -426
rect 199 -498 204 -493
rect 73 -519 78 -514
rect 1933 595 1938 600
rect 972 572 977 577
rect 1804 573 1809 578
rect 846 551 851 556
rect 1611 567 1616 572
rect 1482 545 1487 550
rect 1767 546 1772 551
rect 1638 524 1643 529
rect 1196 507 1201 512
rect 1070 486 1075 491
rect 1769 438 1774 443
rect 1640 416 1645 421
rect 1935 401 1940 406
rect 997 357 1002 362
rect 845 337 850 342
rect 1186 316 1191 321
rect 1034 296 1039 301
rect 975 281 980 286
rect 849 260 854 265
rect 1013 183 1018 188
rect 831 159 836 164
rect 1229 134 1234 139
rect 1052 114 1057 119
rect 993 94 998 99
rect 841 74 846 79
rect 971 29 976 34
rect 845 8 850 13
rect 1806 379 1811 384
rect 1613 373 1618 378
rect 1484 351 1489 356
rect 1769 352 1774 357
rect 1640 330 1645 335
rect 1776 237 1781 242
rect 1647 215 1652 220
rect 1942 200 1947 205
rect 1813 178 1818 183
rect 1620 172 1625 177
rect 1491 150 1496 155
rect 1776 151 1781 156
rect 1647 129 1652 134
rect 980 -331 985 -326
rect 798 -354 803 -349
rect 823 -504 828 -499
rect 834 -640 839 -635
rect 1264 -416 1269 -411
rect 1082 -439 1087 -434
rect 1000 -484 1005 -479
rect 986 -620 991 -615
rect 975 -702 980 -697
rect 849 -723 854 -718
<< metal3 >>
rect -28 1016 132 1017
rect -28 1013 298 1016
rect -28 911 -24 1013
rect -28 906 -26 911
rect 9 732 13 1013
rect 69 871 73 1013
rect 128 1012 298 1013
rect 128 976 132 1012
rect 260 998 264 1002
rect 128 971 130 976
rect 294 941 298 1012
rect 426 961 430 965
rect 294 939 299 941
rect 294 938 296 939
rect 104 933 108 937
rect 128 934 296 938
rect 128 893 132 934
rect 1480 930 1640 931
rect 1480 927 1806 930
rect 260 912 264 916
rect 451 893 494 897
rect 128 890 133 893
rect 128 885 130 890
rect 451 871 455 893
rect 69 867 455 871
rect 69 806 73 867
rect 230 823 234 827
rect 1480 825 1484 927
rect 1480 820 1482 825
rect 69 802 107 806
rect 484 805 492 809
rect 9 728 1027 732
rect 9 666 13 728
rect 1023 722 1027 728
rect 1522 722 1526 927
rect 1636 926 1806 927
rect 1636 890 1640 926
rect 1768 912 1772 916
rect 1636 885 1638 890
rect 1802 855 1806 926
rect 1934 875 1938 879
rect 1802 853 1807 855
rect 1802 852 1804 853
rect 1612 847 1616 851
rect 1636 848 1804 852
rect 1636 807 1640 848
rect 1768 826 1772 830
rect 1636 804 1641 807
rect 1636 799 1638 804
rect 1023 718 1526 722
rect -21 665 139 666
rect -21 662 305 665
rect -21 560 -17 662
rect -21 555 -19 560
rect 9 325 13 662
rect 76 455 80 662
rect 135 661 305 662
rect 135 625 139 661
rect 267 647 271 651
rect 135 620 137 625
rect 301 590 305 661
rect 433 610 437 614
rect 301 588 306 590
rect 301 587 303 588
rect 111 582 115 586
rect 135 583 303 587
rect 135 547 139 583
rect 973 577 977 581
rect 267 561 271 565
rect 838 556 850 560
rect 135 546 150 547
rect 135 543 497 546
rect 135 539 140 543
rect 146 542 497 543
rect 135 534 137 539
rect 838 496 842 556
rect 1023 496 1027 718
rect 1522 656 1526 718
rect 1480 655 1640 656
rect 1480 652 1806 655
rect 1480 550 1484 652
rect 1480 545 1482 550
rect 1197 512 1201 516
rect 838 492 1075 496
rect 237 472 241 476
rect 76 451 114 455
rect 487 454 495 458
rect 841 347 845 492
rect 998 362 1002 366
rect 841 342 849 347
rect -51 324 109 325
rect -51 321 275 324
rect -51 219 -47 321
rect -51 214 -49 219
rect 9 -17 13 321
rect 46 173 50 321
rect 105 320 275 321
rect 105 284 109 320
rect 237 306 241 310
rect 105 279 107 284
rect 271 249 275 320
rect 841 307 845 342
rect 1034 307 1038 492
rect 1061 491 1075 492
rect 1061 490 1070 491
rect 1522 462 1526 652
rect 1636 651 1806 652
rect 1636 615 1640 651
rect 1768 637 1772 641
rect 1636 610 1638 615
rect 1802 580 1806 651
rect 1934 600 1938 604
rect 1802 578 1807 580
rect 1802 577 1804 578
rect 1612 572 1616 576
rect 1636 573 1804 577
rect 1636 532 1640 573
rect 1768 551 1772 555
rect 1636 529 1641 532
rect 1636 524 1638 529
rect 1482 461 1642 462
rect 1482 458 1808 461
rect 1482 356 1486 458
rect 1482 351 1484 356
rect 1187 321 1191 325
rect 841 303 1038 307
rect 403 269 407 273
rect 841 269 845 303
rect 1034 301 1038 303
rect 976 286 980 290
rect 1034 290 1038 296
rect 1034 286 1056 290
rect 841 268 854 269
rect 823 265 854 268
rect 823 264 849 265
rect 271 247 276 249
rect 271 246 273 247
rect 81 241 85 245
rect 105 242 273 246
rect 105 201 109 242
rect 237 220 241 224
rect 419 201 478 205
rect 105 198 110 201
rect 105 193 107 198
rect 419 173 423 201
rect 45 169 423 173
rect 46 114 50 169
rect 823 168 827 264
rect 1014 188 1018 192
rect 823 164 836 168
rect 830 163 831 164
rect 831 155 835 159
rect 831 151 841 155
rect 207 131 211 135
rect 46 110 84 114
rect 469 113 477 117
rect 837 84 841 151
rect 1052 119 1056 286
rect 1522 261 1526 458
rect 1638 457 1808 458
rect 1638 421 1642 457
rect 1770 443 1774 447
rect 1638 416 1640 421
rect 1804 386 1808 457
rect 1936 406 1940 410
rect 1804 384 1809 386
rect 1804 383 1806 384
rect 1614 378 1618 382
rect 1638 379 1806 383
rect 1638 338 1642 379
rect 1770 357 1774 361
rect 1638 335 1643 338
rect 1638 330 1640 335
rect 1489 260 1649 261
rect 1489 257 1815 260
rect 1489 155 1493 257
rect 1645 256 1815 257
rect 1645 220 1649 256
rect 1777 242 1781 246
rect 1645 215 1647 220
rect 1811 185 1815 256
rect 1943 205 1947 209
rect 1811 183 1816 185
rect 1811 182 1813 183
rect 1621 177 1625 181
rect 1645 178 1813 182
rect 1489 150 1491 155
rect 1230 139 1234 143
rect 1645 137 1649 178
rect 1777 156 1781 160
rect 1645 134 1650 137
rect 1645 129 1647 134
rect 994 99 998 103
rect 837 79 845 84
rect 837 74 841 79
rect 842 49 846 74
rect 840 17 846 49
rect 972 34 976 38
rect 840 13 850 17
rect 840 8 845 13
rect 840 5 848 8
rect -52 -18 108 -17
rect -52 -21 274 -18
rect -52 -123 -48 -21
rect -52 -128 -50 -123
rect 9 -299 13 -21
rect 45 -162 49 -21
rect 104 -22 274 -21
rect 104 -58 108 -22
rect 236 -36 240 -32
rect 104 -63 106 -58
rect 270 -93 274 -22
rect 840 -49 844 5
rect 779 -53 844 -49
rect 402 -73 406 -69
rect 270 -95 275 -93
rect 270 -96 272 -95
rect 80 -101 84 -97
rect 104 -100 272 -96
rect 104 -141 108 -100
rect 236 -122 240 -118
rect 446 -141 469 -137
rect 104 -144 109 -141
rect 104 -149 106 -144
rect 446 -162 450 -141
rect 45 -166 450 -162
rect 45 -228 49 -166
rect 206 -211 210 -207
rect 45 -232 83 -228
rect 460 -229 468 -225
rect -58 -300 102 -299
rect -58 -303 268 -300
rect -58 -405 -54 -303
rect -58 -410 -56 -405
rect 39 -510 43 -303
rect 98 -304 268 -303
rect 98 -340 102 -304
rect 230 -318 234 -314
rect 98 -345 100 -340
rect 264 -375 268 -304
rect 779 -341 783 -53
rect 981 -326 985 -322
rect 779 -345 799 -341
rect 396 -355 400 -351
rect 264 -377 269 -375
rect 264 -378 266 -377
rect 74 -383 78 -379
rect 98 -382 266 -378
rect 98 -423 102 -382
rect 230 -404 234 -400
rect 98 -426 103 -423
rect 98 -431 100 -426
rect 779 -430 783 -345
rect 795 -349 803 -345
rect 795 -350 798 -349
rect 1265 -411 1269 -407
rect 1079 -430 1083 -426
rect 779 -434 1087 -430
rect 200 -493 204 -489
rect 39 -514 77 -510
rect 799 -519 803 -434
rect 823 -499 827 -434
rect 1079 -435 1082 -434
rect 1001 -479 1005 -475
rect 799 -523 834 -519
rect 830 -630 834 -523
rect 987 -615 991 -611
rect 830 -631 838 -630
rect 819 -635 838 -631
rect 819 -713 823 -635
rect 830 -640 834 -635
rect 835 -641 839 -640
rect 976 -697 980 -693
rect 819 -717 854 -713
rect 840 -718 854 -717
rect 840 -719 849 -718
<< m4contact >>
rect 259 1002 264 1007
rect 103 937 108 942
rect 425 965 430 970
rect 259 916 264 921
rect 229 827 234 832
rect 479 804 484 809
rect 1767 916 1772 921
rect 1611 851 1616 856
rect 1933 879 1938 884
rect 1767 830 1772 835
rect 266 651 271 656
rect 110 586 115 591
rect 432 614 437 619
rect 972 581 977 586
rect 266 565 271 570
rect 1196 516 1201 521
rect 236 476 241 481
rect 482 453 487 458
rect 997 366 1002 371
rect 236 310 241 315
rect 80 245 85 250
rect 1767 641 1772 646
rect 1611 576 1616 581
rect 1933 604 1938 609
rect 1767 555 1772 560
rect 1186 325 1191 330
rect 402 273 407 278
rect 975 290 980 295
rect 236 224 241 229
rect 1013 192 1018 197
rect 206 135 211 140
rect 464 112 469 117
rect 1769 447 1774 452
rect 1613 382 1618 387
rect 1935 410 1940 415
rect 1769 361 1774 366
rect 1776 246 1781 251
rect 1620 181 1625 186
rect 1942 209 1947 214
rect 1229 143 1234 148
rect 1776 160 1781 165
rect 993 103 998 108
rect 971 38 976 43
rect 235 -32 240 -27
rect 79 -97 84 -92
rect 401 -69 406 -64
rect 235 -118 240 -113
rect 205 -207 210 -202
rect 455 -230 460 -225
rect 229 -314 234 -309
rect 73 -379 78 -374
rect 980 -322 985 -317
rect 395 -351 400 -346
rect 229 -400 234 -395
rect 1264 -407 1269 -402
rect 199 -489 204 -484
rect 1000 -475 1005 -470
rect 986 -611 991 -606
rect 975 -693 980 -688
<< metal4 >>
rect 264 1003 272 1007
rect 268 942 272 1003
rect 430 966 438 970
rect 108 938 272 942
rect 268 921 272 938
rect 264 920 272 921
rect 434 920 438 966
rect 264 917 438 920
rect 268 916 438 917
rect 1772 917 1780 921
rect 281 832 285 916
rect 234 828 285 832
rect 345 807 349 916
rect 1776 856 1780 917
rect 1938 880 1946 884
rect 1616 852 1780 856
rect 1776 835 1780 852
rect 1772 834 1780 835
rect 1942 834 1946 880
rect 1772 831 1946 834
rect 1776 830 1946 831
rect 477 807 479 809
rect 345 804 479 807
rect 345 803 481 804
rect 345 697 349 803
rect 345 693 1077 697
rect 271 652 279 656
rect 275 591 279 652
rect 115 587 279 591
rect 275 570 279 587
rect 271 569 279 570
rect 345 569 349 693
rect 1073 685 1077 693
rect 1876 685 1880 830
rect 1073 681 1880 685
rect 437 615 445 619
rect 441 569 445 615
rect 1073 586 1077 681
rect 1772 642 1780 646
rect 977 582 1208 586
rect 271 566 445 569
rect 275 565 445 566
rect 288 481 292 565
rect 241 477 292 481
rect 345 458 349 565
rect 345 453 482 458
rect 241 311 249 315
rect 245 250 249 311
rect 85 246 249 250
rect 245 229 249 246
rect 241 228 249 229
rect 345 228 349 453
rect 1005 371 1009 582
rect 1204 521 1208 582
rect 1776 581 1780 642
rect 1616 577 1780 581
rect 1776 560 1780 577
rect 1772 559 1780 560
rect 1876 559 1880 681
rect 1938 605 1946 609
rect 1942 559 1946 605
rect 1772 556 1946 559
rect 1776 555 1946 556
rect 1201 517 1208 521
rect 1205 513 1241 517
rect 1002 368 1010 371
rect 1002 367 1198 368
rect 1006 364 1198 367
rect 1018 295 1022 364
rect 1194 330 1198 364
rect 1191 326 1198 330
rect 980 291 1025 295
rect 407 274 415 278
rect 411 228 415 274
rect 241 225 415 228
rect 245 224 415 225
rect 258 140 262 224
rect 211 136 262 140
rect 345 117 349 224
rect 1021 197 1025 291
rect 1018 193 1025 197
rect 1022 188 1025 193
rect 345 113 464 117
rect 240 -31 248 -27
rect 244 -92 248 -31
rect 84 -96 248 -92
rect 244 -113 248 -96
rect 240 -114 248 -113
rect 345 -114 349 113
rect 1021 108 1025 188
rect 1237 148 1241 513
rect 1774 448 1782 452
rect 1778 387 1782 448
rect 1618 383 1782 387
rect 1778 366 1782 383
rect 1774 365 1782 366
rect 1876 365 1880 555
rect 1940 411 1948 415
rect 1944 365 1948 411
rect 1774 362 1948 365
rect 1778 361 1948 362
rect 1781 247 1789 251
rect 1785 186 1789 247
rect 1625 182 1789 186
rect 1785 165 1789 182
rect 1781 164 1789 165
rect 1876 164 1880 361
rect 1947 210 1955 214
rect 1951 164 1955 210
rect 1781 161 1955 164
rect 1785 160 1955 161
rect 1234 144 1241 148
rect 998 104 1025 108
rect 1016 43 1020 104
rect 976 41 1020 43
rect 976 39 1200 41
rect 1014 37 1200 39
rect 406 -68 414 -64
rect 410 -114 414 -68
rect 240 -117 414 -114
rect 244 -118 414 -117
rect 257 -202 261 -118
rect 210 -206 261 -202
rect 345 -225 349 -118
rect 345 -229 455 -225
rect 234 -313 242 -309
rect 238 -374 242 -313
rect 78 -378 242 -374
rect 238 -395 242 -378
rect 234 -396 242 -395
rect 345 -396 349 -229
rect 1196 -317 1200 37
rect 985 -321 1292 -317
rect 400 -350 408 -346
rect 404 -396 408 -350
rect 234 -399 408 -396
rect 238 -400 408 -399
rect 251 -484 255 -400
rect 1008 -461 1012 -321
rect 1269 -403 1273 -402
rect 1288 -403 1292 -321
rect 1269 -406 1292 -403
rect 1277 -407 1292 -406
rect 1008 -465 1026 -461
rect 1008 -470 1012 -465
rect 1005 -474 1012 -470
rect 204 -488 255 -484
rect 1022 -506 1026 -465
rect 993 -510 1026 -506
rect 993 -600 997 -510
rect 993 -604 1010 -600
rect 993 -606 997 -604
rect 991 -610 997 -606
rect 1006 -675 1010 -604
rect 983 -679 1010 -675
rect 983 -688 987 -679
rect 980 -692 987 -688
<< labels >>
rlabel metal1 -72 931 -68 935 1 a0
rlabel metal1 -72 913 -68 917 1 b0
rlabel metal1 -65 580 -61 584 1 a1
rlabel metal1 -65 562 -61 566 1 b1
rlabel metal1 -95 239 -91 243 1 a2
rlabel metal1 -95 221 -91 225 1 b2
rlabel metal1 -96 -103 -92 -99 1 a3
rlabel metal1 -96 -121 -92 -117 1 b3
rlabel metal1 -102 -385 -98 -381 3 a4
rlabel metal1 -102 -403 -98 -399 3 b4
rlabel metal1 479 836 483 840 1 gn0
rlabel metal1 484 626 488 630 7 p1
rlabel metal1 486 485 490 489 7 gn1
rlabel metal1 454 285 458 289 1 p2
rlabel metal1 456 144 460 148 1 gn2
rlabel metal1 453 -57 457 -53 1 p3
rlabel metal1 455 -198 459 -194 1 gn3
rlabel metal1 447 -339 451 -335 1 p4
rlabel metal1 449 -480 453 -476 1 gn4
rlabel metal1 534 836 538 840 7 g0
rlabel metal1 537 485 541 489 7 g1
rlabel metal1 516 144 520 148 1 g2
rlabel metal1 510 -198 514 -194 1 g3
rlabel metal1 1390 193 1394 197 1 c4
rlabel metal1 1386 379 1390 383 1 c3
rlabel metal1 1384 538 1388 542 1 c2
rlabel metal1 477 977 481 981 1 s0
rlabel metal1 1377 835 1381 839 1 c1
rlabel metal3 43 1013 47 1017 5 vdd
rlabel metal4 434 929 438 933 1 gnd
rlabel metal1 1875 888 1879 892 1 s1
rlabel metal1 1875 613 1879 617 1 s2
rlabel metal1 1877 419 1881 423 1 s3
rlabel metal1 1884 218 1888 222 1 s4
rlabel metal1 1480 -361 1484 -357 1 cout
<< end >>
