magic
tech scmos
timestamp 1763399017
<< nwell >>
rect 10 -34 43 59
rect 62 -20 88 32
rect 122 -20 148 32
rect 182 -34 206 18
<< ntransistor >>
rect 21 -83 23 -63
rect 73 -69 75 -29
rect 81 -69 83 -29
rect 133 -69 135 -29
rect 141 -69 143 -29
rect 193 -62 195 -42
<< ptransistor >>
rect 21 -27 23 53
rect 29 -27 31 53
rect 73 -14 75 26
rect 133 -14 135 26
rect 193 -28 195 12
<< ndiffusion >>
rect 20 -83 21 -63
rect 23 -83 24 -63
rect 28 -83 29 -63
rect 72 -69 73 -29
rect 75 -69 76 -29
rect 80 -69 81 -29
rect 83 -69 84 -29
rect 132 -69 133 -29
rect 135 -69 136 -29
rect 140 -69 141 -29
rect 143 -69 144 -29
rect 192 -62 193 -42
rect 195 -62 196 -42
<< pdiffusion >>
rect 20 -27 21 53
rect 23 -27 24 53
rect 28 -27 29 53
rect 31 -27 32 53
rect 36 -27 37 53
rect 72 -14 73 26
rect 75 -14 76 26
rect 132 -14 133 26
rect 135 -14 136 26
rect 192 -28 193 12
rect 195 -28 196 12
<< ndcontact >>
rect 16 -83 20 -63
rect 24 -83 28 -63
rect 68 -69 72 -29
rect 76 -69 80 -29
rect 84 -69 88 -29
rect 128 -69 132 -29
rect 136 -69 140 -29
rect 144 -69 148 -29
rect 188 -62 192 -42
rect 196 -62 200 -42
<< pdcontact >>
rect 16 -27 20 53
rect 24 -27 28 53
rect 32 -27 36 53
rect 68 -14 72 26
rect 76 -14 80 26
rect 128 -14 132 26
rect 136 -14 140 26
rect 188 -28 192 12
rect 196 -28 200 12
<< polysilicon >>
rect 21 53 23 66
rect 29 53 31 66
rect 73 26 75 37
rect 133 26 135 37
rect 193 12 195 15
rect 21 -63 23 -27
rect 29 -38 31 -27
rect 73 -29 75 -14
rect 81 -29 83 -26
rect 133 -29 135 -14
rect 141 -29 143 -26
rect 193 -42 195 -28
rect 193 -65 195 -62
rect 73 -73 75 -69
rect 81 -73 83 -69
rect 133 -73 135 -69
rect 141 -73 143 -69
rect 21 -93 23 -83
<< polycontact >>
rect 20 66 24 70
rect 28 66 32 70
rect 72 37 76 41
rect 132 37 136 41
rect 80 -26 84 -22
rect 140 -26 144 -22
rect 189 -39 193 -35
<< metal1 >>
rect -10 89 187 95
rect -10 53 -4 89
rect 4 78 62 83
rect 4 58 9 78
rect 20 70 24 73
rect 28 70 76 73
rect 4 53 20 58
rect -11 47 8 53
rect -12 23 1 29
rect -4 -86 1 23
rect 24 53 28 58
rect 72 46 76 70
rect 72 41 113 46
rect 62 32 67 36
rect 62 27 72 32
rect 67 26 72 27
rect 67 23 68 26
rect 101 -10 105 -5
rect 80 -14 105 -10
rect 51 -26 80 -22
rect 32 -41 38 -27
rect 51 -41 58 -26
rect 101 -29 105 -14
rect 108 -21 113 41
rect 119 29 125 89
rect 119 26 131 29
rect 119 23 128 26
rect 181 20 187 89
rect 181 16 206 20
rect 188 12 192 16
rect 136 -17 175 -14
rect 108 -22 142 -21
rect 108 -26 140 -22
rect 24 -44 58 -41
rect 24 -47 57 -44
rect 24 -63 29 -47
rect 66 -79 71 -69
rect 76 -74 80 -69
rect 101 -69 107 -29
rect 84 -73 107 -69
rect 16 -86 20 -83
rect 66 -84 74 -79
rect -4 -91 20 -86
rect 14 -104 19 -91
rect 69 -103 74 -84
rect 127 -103 132 -69
rect 136 -74 140 -69
rect 171 -36 178 -17
rect 182 -36 189 -35
rect 165 -39 189 -36
rect 196 -36 200 -28
rect 165 -41 182 -39
rect 196 -40 206 -36
rect 144 -81 149 -69
rect 165 -81 170 -41
rect 196 -42 200 -40
rect 188 -71 192 -62
rect 182 -75 206 -71
rect 144 -86 170 -81
rect 183 -103 188 -75
rect 69 -104 188 -103
rect 14 -108 188 -104
rect 14 -109 74 -108
<< m2contact >>
rect 62 78 67 83
rect 62 36 67 41
rect 100 -5 105 0
rect 132 41 137 46
<< metal2 >>
rect 62 41 67 78
rect 101 41 132 45
rect 101 0 105 41
<< labels >>
rlabel metal1 -11 47 -3 53 3 vdd
rlabel metal1 -12 23 -4 29 3 gnd
rlabel metal1 40 70 55 72 1 clk
rlabel metal1 200 -40 205 -36 7 q
rlabel metal1 20 70 23 72 1 d
rlabel metal1 172 -36 176 -20 1 q_int
rlabel metal1 54 -44 58 -28 1 x1
rlabel metal1 24 53 28 58 1 x2
rlabel metal1 103 -45 107 -40 1 y
rlabel metal1 76 -74 80 -69 1 x3
rlabel metal1 136 -74 140 -69 1 x4
rlabel metal1 10 54 14 56 1 vdd
rlabel metal1 183 44 185 71 1 vdd
rlabel metal1 6 92 155 93 5 vdd
rlabel metal2 62 47 65 51 1 vdd
<< end >>
