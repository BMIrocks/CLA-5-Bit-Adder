**5-bit Carry Lookahead Adder Block
.include INV.cir
.include NAND2.cir
.include XOR2.cir
.include PG.cir
.include CARRY.cir

.subckt CLA a0 a1 a2 a3 a4 b0 b1 b2 b3 b4 s0 s1 s2 s3 s4 cout vdd gnd
* Propagate and Generate
XPG0 a0 b0 p0 g0n vdd gnd PG
XPG1 a1 b1 p1 g1n vdd gnd PG
XPG2 a2 b2 p2 g2n vdd gnd PG
XPG3 a3 b3 p3 g3n vdd gnd PG
XPG4 a4 b4 p4 g4n vdd gnd PG

* Carry
XCARRY p0 p1 p2 p3 p4 g0n g1n g2n g3n g4n c1 c2 c3 c4 cout vdd gnd CARRY

* Sum
XXOR0 p0 gnd s0 vdd gnd XOR2
XXOR1 p1 c1 s1 vdd gnd XOR2
XXOR2 p2 c2 s2 vdd gnd XOR2
XXOR3 p3 c3 s3 vdd gnd XOR2
XXOR4 p4 c4 s4 vdd gnd XOR2
.ends CLA